
module cht ( v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, 
        f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, 
        j, i, h, g, f, e, d, c, a, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, 
        u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, 
        c1, b1, a1, z0, y0, x0, w0 );
  input v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0,
         d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i,
         h, g, f, e, d, c, a;
  output f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1,
         o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0,
         x0, w0;
  wire   n6, n7, n8, n9, n12, n13, n23, n24, n25, n26, n27, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n67, n68, n71, n72, n75, n76, n79, n80, n81, n84, n85,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150;

  or2 U4 ( .A1(n6), .A2(n7), .Z(z0) );
  and2 U5 ( .A1(c), .A2(n8), .Z(n7) );
  and2 U6 ( .A1(p), .A2(n9), .Z(n6) );
  or2 U10 ( .A1(n12), .A2(n13), .Z(y0) );
  and2 U11 ( .A1(h), .A2(n8), .Z(n13) );
  and2 U12 ( .A1(o), .A2(n9), .Z(n12) );
  or2 U20 ( .A1(n23), .A2(n24), .Z(x0) );
  and2 U21 ( .A1(g), .A2(n8), .Z(n24) );
  and2 U22 ( .A1(n), .A2(n9), .Z(n23) );
  or2 U23 ( .A1(n25), .A2(n26), .Z(w1) );
  and2 U24 ( .A1(n27), .A2(n0), .Z(n26) );
  or2 U26 ( .A1(n29), .A2(n30), .Z(w0) );
  and2 U27 ( .A1(f), .A2(n8), .Z(n30) );
  and2 U28 ( .A1(m), .A2(n9), .Z(n29) );
  or2 U29 ( .A1(n31), .A2(n32), .Z(v1) );
  and2 U30 ( .A1(n27), .A2(m0), .Z(n32) );
  or2 U32 ( .A1(n33), .A2(n34), .Z(u1) );
  and2 U33 ( .A1(l0), .A2(n27), .Z(n34) );
  or2 U35 ( .A1(n35), .A2(n36), .Z(t1) );
  and2 U36 ( .A1(k0), .A2(n27), .Z(n36) );
  or2 U38 ( .A1(n37), .A2(n38), .Z(s1) );
  and2 U39 ( .A1(j0), .A2(n27), .Z(n38) );
  or2 U41 ( .A1(n39), .A2(n40), .Z(r1) );
  and2 U42 ( .A1(i0), .A2(n27), .Z(n40) );
  or2 U44 ( .A1(n41), .A2(n42), .Z(q1) );
  and2 U45 ( .A1(h0), .A2(n27), .Z(n42) );
  or2 U49 ( .A1(n43), .A2(n44), .Z(p1) );
  and2 U50 ( .A1(n45), .A2(a), .Z(n44) );
  and2 U51 ( .A1(f0), .A2(n142), .Z(n43) );
  or2 U52 ( .A1(n47), .A2(n48), .Z(o1) );
  and2 U53 ( .A1(n45), .A2(f0), .Z(n48) );
  and2 U54 ( .A1(e0), .A2(n141), .Z(n47) );
  or2 U55 ( .A1(n49), .A2(n50), .Z(n1) );
  and2 U56 ( .A1(e0), .A2(n145), .Z(n50) );
  and2 U57 ( .A1(d0), .A2(n142), .Z(n49) );
  or2 U58 ( .A1(n51), .A2(n52), .Z(m1) );
  and2 U59 ( .A1(d0), .A2(n145), .Z(n52) );
  and2 U60 ( .A1(c0), .A2(n143), .Z(n51) );
  or2 U61 ( .A1(n53), .A2(n54), .Z(l1) );
  and2 U62 ( .A1(c0), .A2(n45), .Z(n54) );
  and2 U63 ( .A1(b0), .A2(n142), .Z(n53) );
  or2 U64 ( .A1(n55), .A2(n56), .Z(k1) );
  and2 U65 ( .A1(b0), .A2(n145), .Z(n56) );
  and2 U66 ( .A1(a0), .A2(n143), .Z(n55) );
  or2 U67 ( .A1(n57), .A2(n58), .Z(j1) );
  and2 U68 ( .A1(a0), .A2(n45), .Z(n58) );
  and2 U69 ( .A1(z), .A2(n142), .Z(n57) );
  or2 U70 ( .A1(n59), .A2(n60), .Z(i1) );
  and2 U71 ( .A1(z), .A2(n145), .Z(n60) );
  and2 U72 ( .A1(y), .A2(n143), .Z(n59) );
  or2 U73 ( .A1(n61), .A2(n62), .Z(h1) );
  and2 U74 ( .A1(y), .A2(n145), .Z(n62) );
  and2 U75 ( .A1(x), .A2(n142), .Z(n61) );
  or2 U76 ( .A1(n63), .A2(n64), .Z(g1) );
  and2 U77 ( .A1(x), .A2(n45), .Z(n64) );
  and2 U78 ( .A1(w), .A2(n141), .Z(n63) );
  or2 U82 ( .A1(n67), .A2(n68), .Z(f1) );
  and2 U83 ( .A1(w), .A2(n45), .Z(n68) );
  and2 U84 ( .A1(v), .A2(n141), .Z(n67) );
  or2 U88 ( .A1(n71), .A2(n72), .Z(e1) );
  and2 U89 ( .A1(v), .A2(n45), .Z(n72) );
  and2 U90 ( .A1(u), .A2(n141), .Z(n71) );
  or2 U94 ( .A1(n75), .A2(n76), .Z(d1) );
  and2 U95 ( .A1(u), .A2(n45), .Z(n76) );
  and2 U96 ( .A1(t), .A2(n141), .Z(n75) );
  or2 U100 ( .A1(n79), .A2(n80), .Z(c1) );
  and2 U101 ( .A1(t), .A2(n45), .Z(n80) );
  and2 U103 ( .A1(s), .A2(n143), .Z(n79) );
  or2 U109 ( .A1(n84), .A2(n85), .Z(b1) );
  and2 U110 ( .A1(e), .A2(n8), .Z(n85) );
  and2 U111 ( .A1(r), .A2(n9), .Z(n84) );
  or2 U120 ( .A1(n89), .A2(n90), .Z(a1) );
  and2 U121 ( .A1(d), .A2(n8), .Z(n90) );
  and2 U122 ( .A1(n140), .A2(i), .Z(n8) );
  and2 U123 ( .A1(q), .A2(n9), .Z(n89) );
  and2 U124 ( .A1(n140), .A2(n91), .Z(n9) );
  inv1 U125 ( .I(i), .ZN(n91) );
  inv1 U128 ( .I(n92), .ZN(n45) );
  inv1 U129 ( .I(n110), .ZN(n93) );
  inv1 U132 ( .I(g0), .ZN(n94) );
  or2 U133 ( .A1(n113), .A2(n94), .Z(n95) );
  inv1 U134 ( .I(n95), .ZN(n41) );
  inv1 U135 ( .I(h0), .ZN(n96) );
  or2 U136 ( .A1(n113), .A2(n96), .Z(n97) );
  inv1 U137 ( .I(n97), .ZN(n39) );
  inv1 U138 ( .I(i0), .ZN(n98) );
  or2 U139 ( .A1(n113), .A2(n98), .Z(n99) );
  inv1 U140 ( .I(n99), .ZN(n37) );
  inv1 U141 ( .I(j0), .ZN(n100) );
  or2 U142 ( .A1(n113), .A2(n100), .Z(n101) );
  inv1 U143 ( .I(n101), .ZN(n35) );
  inv1 U144 ( .I(k0), .ZN(n102) );
  or2 U145 ( .A1(n113), .A2(n102), .Z(n103) );
  inv1 U146 ( .I(n103), .ZN(n33) );
  inv1 U147 ( .I(l0), .ZN(n104) );
  or2 U148 ( .A1(n113), .A2(n104), .Z(n105) );
  inv1 U149 ( .I(n105), .ZN(n31) );
  inv1 U150 ( .I(m0), .ZN(n106) );
  or2 U151 ( .A1(n113), .A2(n106), .Z(n107) );
  inv1 U152 ( .I(n107), .ZN(n25) );
  and2 U157 ( .A1(o0), .A2(n93), .Z(n118) );
  and2 U158 ( .A1(p), .A2(k), .Z(n112) );
  and2 U159 ( .A1(a), .A2(n140), .Z(n111) );
  and2 U160 ( .A1(n112), .A2(n111), .Z(n116) );
  and2 U162 ( .A1(n147), .A2(n0), .Z(n115) );
  or2 U164 ( .A1(n118), .A2(n117), .Z(x1) );
  inv1 U165 ( .I(p), .ZN(n119) );
  and2 U169 ( .A1(o0), .A2(n146), .Z(n123) );
  and2 U170 ( .A1(p0), .A2(n93), .Z(n122) );
  or2 U171 ( .A1(n123), .A2(n122), .Z(y1) );
  and2 U172 ( .A1(p0), .A2(n146), .Z(n125) );
  and2 U173 ( .A1(q0), .A2(n150), .Z(n124) );
  or2 U174 ( .A1(n125), .A2(n124), .Z(z1) );
  and2 U175 ( .A1(q0), .A2(n146), .Z(n127) );
  and2 U176 ( .A1(r0), .A2(n137), .Z(n126) );
  or2 U177 ( .A1(n127), .A2(n126), .Z(a2) );
  and2 U178 ( .A1(r0), .A2(n146), .Z(n129) );
  and2 U179 ( .A1(s0), .A2(n137), .Z(n128) );
  or2 U180 ( .A1(n129), .A2(n128), .Z(b2) );
  and2 U181 ( .A1(s0), .A2(n146), .Z(n131) );
  and2 U182 ( .A1(t0), .A2(n150), .Z(n130) );
  or2 U183 ( .A1(n131), .A2(n130), .Z(c2) );
  and2 U184 ( .A1(t0), .A2(n146), .Z(n133) );
  and2 U185 ( .A1(u0), .A2(n150), .Z(n132) );
  or2 U186 ( .A1(n133), .A2(n132), .Z(d2) );
  and2 U187 ( .A1(u0), .A2(n146), .Z(n135) );
  and2 U188 ( .A1(v0), .A2(n93), .Z(n134) );
  or2 U189 ( .A1(n135), .A2(n134), .Z(e2) );
  and2 U190 ( .A1(v0), .A2(n146), .Z(n139) );
  and2 U191 ( .A1(a), .A2(n137), .Z(n138) );
  or2 U192 ( .A1(n139), .A2(n138), .Z(f2) );
  and2f U127 ( .A1(n140), .A2(k), .Z(n27) );
  or2 U130 ( .A1(l), .A2(j), .Z(n149) );
  inv1 U131 ( .I(n149), .ZN(n141) );
  inv1 U153 ( .I(n149), .ZN(n143) );
  inv1 U154 ( .I(n149), .ZN(n142) );
  inv1 U155 ( .I(j), .ZN(n81) );
  inv1 U156 ( .I(l), .ZN(n148) );
  and2f U161 ( .A1(n119), .A2(k), .Z(n120) );
  or2f U163 ( .A1(n116), .A2(n115), .Z(n117) );
  or2f U166 ( .A1(n109), .A2(p), .Z(n144) );
  or2f U167 ( .A1(l), .A2(n108), .Z(n109) );
  inv1 U168 ( .I(n92), .ZN(n145) );
  or2f U193 ( .A1(l), .A2(n81), .Z(n92) );
  inv1f U194 ( .I(n121), .ZN(n146) );
  or2f U195 ( .A1(n120), .A2(l), .Z(n121) );
  and2f U196 ( .A1(n148), .A2(n108), .Z(n147) );
  inv1 U197 ( .I(n147), .ZN(n113) );
  inv1f U198 ( .I(k), .ZN(n108) );
  inv1f U199 ( .I(l), .ZN(n140) );
  inv1f U200 ( .I(n144), .ZN(n150) );
  inv1f U201 ( .I(n144), .ZN(n137) );
  or2f U202 ( .A1(n109), .A2(p), .Z(n110) );
endmodule

