
module i8 ( V118, V122, V119, V121, V51, V52, V50, V116, V49, V48, V15, V84, 
        V47, V133, V214, V213, V212, V197, V165, V150, V149, V146, V145, V143, 
        V142, V136, V134 );
  input [1:0] V118;
  input [0:0] V122;
  input [0:0] V119;
  input [17:16] V121;
  input [0:0] V51;
  input [0:0] V52;
  input [0:0] V50;
  input [31:0] V116;
  input [0:0] V49;
  input [0:0] V48;
  input [14:0] V15;
  input [31:0] V84;
  input [31:0] V47;
  input [10:0] V133;
  output [0:0] V214;
  output [0:0] V213;
  output [14:0] V212;
  output [31:0] V197;
  output [14:0] V165;
  output [0:0] V150;
  output [2:0] V149;
  output [0:0] V146;
  output [1:0] V145;
  output [0:0] V143;
  output [5:0] V142;
  output [1:0] V136;
  output [0:0] V134;
  wire   n1, n2, n7, n10, n11, n12, n20, n21, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n68, n71, n72, n73,
         n77, n382, n386, n392, n395, n396, n630, n631, n752, n758, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n771, n772, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n789, n790, n791, n792, n794, n795, n796, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n809, n810, n811, n812,
         n813, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n832, n834, n835, n836, n837, n842, n843, n844, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n874, n875, n876, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753;

  or2 U1 ( .A1(n1), .A2(n2), .Z(V214[0]) );
  and2 U6 ( .A1(V133[10]), .A2(V122[0]), .Z(n7) );
  or2 U8 ( .A1(n10), .A2(n11), .Z(V213[0]) );
  and2 U9 ( .A1(V121[16]), .A2(n12), .Z(n11) );
  or2 U16 ( .A1(n20), .A2(n21), .Z(V212[9]) );
  or2 U17 ( .A1(n858), .A2(n23), .Z(n21) );
  and2 U18 ( .A1(V84[26]), .A2(n24), .Z(n20) );
  or2 U19 ( .A1(n25), .A2(n26), .Z(V212[8]) );
  or2 U20 ( .A1(n858), .A2(n27), .Z(n26) );
  and2 U21 ( .A1(V84[25]), .A2(n24), .Z(n25) );
  or2 U22 ( .A1(n28), .A2(n29), .Z(V212[7]) );
  or2 U23 ( .A1(n858), .A2(n30), .Z(n29) );
  and2 U24 ( .A1(V84[24]), .A2(n24), .Z(n28) );
  or2 U25 ( .A1(n31), .A2(n32), .Z(V212[6]) );
  or2 U26 ( .A1(n858), .A2(n33), .Z(n32) );
  and2 U27 ( .A1(V84[23]), .A2(n24), .Z(n31) );
  or2 U28 ( .A1(n34), .A2(n35), .Z(V212[5]) );
  or2 U29 ( .A1(n858), .A2(n36), .Z(n35) );
  and2 U30 ( .A1(V84[22]), .A2(n24), .Z(n34) );
  or2 U31 ( .A1(n37), .A2(n38), .Z(V212[4]) );
  or2 U32 ( .A1(n858), .A2(n39), .Z(n38) );
  and2 U33 ( .A1(V84[21]), .A2(n24), .Z(n37) );
  or2 U34 ( .A1(n40), .A2(n41), .Z(V212[3]) );
  or2 U35 ( .A1(n858), .A2(n42), .Z(n41) );
  and2 U36 ( .A1(V84[20]), .A2(n24), .Z(n40) );
  or2 U37 ( .A1(n43), .A2(n44), .Z(V212[2]) );
  or2 U38 ( .A1(n858), .A2(n45), .Z(n44) );
  and2 U39 ( .A1(V84[19]), .A2(n24), .Z(n43) );
  or2 U40 ( .A1(n46), .A2(n47), .Z(V212[1]) );
  or2 U41 ( .A1(n858), .A2(n48), .Z(n47) );
  and2 U42 ( .A1(V84[18]), .A2(n24), .Z(n46) );
  or2 U43 ( .A1(n49), .A2(n50), .Z(V212[14]) );
  or2 U44 ( .A1(n858), .A2(n51), .Z(n50) );
  and2 U45 ( .A1(V84[31]), .A2(n24), .Z(n49) );
  or2 U46 ( .A1(n52), .A2(n53), .Z(V212[13]) );
  or2 U47 ( .A1(n858), .A2(n54), .Z(n53) );
  and2 U48 ( .A1(V84[30]), .A2(n24), .Z(n52) );
  or2 U49 ( .A1(n55), .A2(n56), .Z(V212[12]) );
  or2 U50 ( .A1(n858), .A2(n57), .Z(n56) );
  and2 U51 ( .A1(V84[29]), .A2(n24), .Z(n55) );
  or2 U52 ( .A1(n58), .A2(n59), .Z(V212[11]) );
  or2 U53 ( .A1(n858), .A2(n60), .Z(n59) );
  and2 U54 ( .A1(V84[28]), .A2(n24), .Z(n58) );
  or2 U55 ( .A1(n61), .A2(n62), .Z(V212[10]) );
  or2 U56 ( .A1(n858), .A2(n63), .Z(n62) );
  and2 U57 ( .A1(V84[27]), .A2(n24), .Z(n61) );
  or2 U58 ( .A1(n64), .A2(n65), .Z(V212[0]) );
  or2 U59 ( .A1(n858), .A2(n66), .Z(n65) );
  or2 U63 ( .A1(V118[0]), .A2(n72), .Z(n71) );
  or2 U64 ( .A1(V118[1]), .A2(n73), .Z(n68) );
  or2 U65 ( .A1(V133[2]), .A2(V133[1]), .Z(n73) );
  and2 U66 ( .A1(V84[17]), .A2(n24), .Z(n64) );
  and2 U374 ( .A1(n386), .A2(n392), .Z(n382) );
  inv1 U375 ( .I(V118[0]), .ZN(n392) );
  or2 U379 ( .A1(V133[10]), .A2(n77), .Z(n395) );
  inv1 U651 ( .I(n631), .ZN(n630) );
  or2 U652 ( .A1(V133[7]), .A2(V133[3]), .Z(n631) );
  and2 U814 ( .A1(n396), .A2(n1739), .Z(n752) );
  or2 U829 ( .A1(V133[9]), .A2(V133[10]), .Z(n758) );
  or2 U833 ( .A1(n761), .A2(n762), .Z(V134[0]) );
  and2 U834 ( .A1(V48[0]), .A2(n763), .Z(n762) );
  and2 U835 ( .A1(n764), .A2(n765), .Z(n761) );
  or2 U836 ( .A1(n766), .A2(n767), .Z(n765) );
  and2 U837 ( .A1(V49[0]), .A2(n760), .Z(n767) );
  inv1 U838 ( .I(n72), .ZN(n760) );
  and2 U839 ( .A1(n768), .A2(n72), .Z(n766) );
  or2 U840 ( .A1(V133[10]), .A2(n769), .Z(n72) );
  or2 U841 ( .A1(V133[9]), .A2(V133[7]), .Z(n769) );
  and2 U843 ( .A1(V84[0]), .A2(V133[10]), .Z(n771) );
  or2 U845 ( .A1(V116[0]), .A2(n1738), .Z(n772) );
  inv1 U858 ( .I(V133[9]), .ZN(n777) );
  and2 U860 ( .A1(n1063), .A2(n1140), .Z(n779) );
  inv1 U864 ( .I(n1024), .ZN(n782) );
  and2 U865 ( .A1(n1403), .A2(n1402), .Z(n783) );
  inv1 U866 ( .I(n783), .ZN(n826) );
  and2 U867 ( .A1(n1600), .A2(n1599), .Z(n784) );
  inv1 U868 ( .I(n784), .ZN(n823) );
  or2 U869 ( .A1(n825), .A2(V133[10]), .Z(n785) );
  and2 U872 ( .A1(n791), .A2(V47[7]), .Z(n787) );
  and2 U874 ( .A1(n791), .A2(V47[9]), .Z(n789) );
  and2 U875 ( .A1(n791), .A2(V47[10]), .Z(n790) );
  inv1 U876 ( .I(n862), .ZN(n791) );
  and2 U877 ( .A1(n799), .A2(V47[11]), .Z(n792) );
  and2 U879 ( .A1(n791), .A2(V47[12]), .Z(n794) );
  and2 U880 ( .A1(n791), .A2(V47[13]), .Z(n795) );
  and2 U881 ( .A1(n799), .A2(V47[14]), .Z(n796) );
  and2 U883 ( .A1(n799), .A2(V47[16]), .Z(n798) );
  inv1 U884 ( .I(n863), .ZN(n799) );
  inv1 U886 ( .I(n800), .ZN(n801) );
  and2 U894 ( .A1(n837), .A2(V84[14]), .Z(n809) );
  and2 U895 ( .A1(n874), .A2(V84[1]), .Z(n810) );
  or2 U896 ( .A1(n1558), .A2(n811), .Z(n1560) );
  or2 U897 ( .A1(n882), .A2(n1559), .Z(n811) );
  or2 U898 ( .A1(n1594), .A2(n812), .Z(n1596) );
  or2 U899 ( .A1(n882), .A2(n1595), .Z(n812) );
  or2 U907 ( .A1(n821), .A2(n822), .Z(n820) );
  inv1 U909 ( .I(n1504), .ZN(n822) );
  or2 U912 ( .A1(n828), .A2(n829), .Z(n827) );
  inv1 U913 ( .I(n1434), .ZN(n828) );
  inv1 U914 ( .I(n1433), .ZN(n829) );
  and2 U915 ( .A1(n837), .A2(V84[11]), .Z(n830) );
  inv1 U919 ( .I(n834), .ZN(n1102) );
  inv1 U921 ( .I(n1034), .ZN(n836) );
  or2 U931 ( .A1(n847), .A2(n848), .Z(n846) );
  inv1 U932 ( .I(n1474), .ZN(n847) );
  inv1 U933 ( .I(n1473), .ZN(n848) );
  or2 U934 ( .A1(n850), .A2(n851), .Z(n849) );
  inv1 U935 ( .I(n1531), .ZN(n850) );
  inv1 U936 ( .I(n1530), .ZN(n851) );
  or2 U937 ( .A1(n825), .A2(n1072), .Z(n852) );
  inv1 U942 ( .I(n786), .ZN(n856) );
  inv1 U945 ( .I(n891), .ZN(n858) );
  inv1 U946 ( .I(n1091), .ZN(n859) );
  inv1 U947 ( .I(n1091), .ZN(n860) );
  inv1 U949 ( .I(n861), .ZN(n862) );
  inv1 U956 ( .I(n868), .ZN(n869) );
  inv1 U959 ( .I(n1529), .ZN(n872) );
  inv1 U963 ( .I(n1358), .ZN(n876) );
  inv1 U968 ( .I(n1362), .ZN(n881) );
  inv1 U969 ( .I(n1362), .ZN(n882) );
  inv1 U970 ( .I(n1362), .ZN(n883) );
  inv1 U972 ( .I(V133[10]), .ZN(n922) );
  and2 U973 ( .A1(n772), .A2(n922), .Z(n884) );
  or2 U974 ( .A1(n884), .A2(n771), .Z(n768) );
  and2 U975 ( .A1(n396), .A2(n922), .Z(n930) );
  or2 U977 ( .A1(n824), .A2(n853), .Z(n981) );
  and2 U978 ( .A1(n930), .A2(n981), .Z(n763) );
  inv1 U979 ( .I(n763), .ZN(n764) );
  inv1 U980 ( .I(V133[8]), .ZN(n1739) );
  inv1 U981 ( .I(n77), .ZN(n885) );
  or2 U985 ( .A1(n1088), .A2(V133[5]), .Z(n1346) );
  and2 U986 ( .A1(n885), .A2(n1346), .Z(n886) );
  or2 U987 ( .A1(n886), .A2(V133[2]), .Z(n887) );
  inv1 U988 ( .I(n887), .ZN(n888) );
  or2 U989 ( .A1(n888), .A2(V133[10]), .Z(n24) );
  inv1 U990 ( .I(V133[5]), .ZN(n889) );
  or2 U991 ( .A1(n889), .A2(n68), .Z(n890) );
  or2 U992 ( .A1(n890), .A2(n71), .Z(n891) );
  or2 U993 ( .A1(n1738), .A2(V133[10]), .Z(n1529) );
  inv1 U994 ( .I(V116[0]), .ZN(n892) );
  or2 U995 ( .A1(n1529), .A2(n892), .Z(n893) );
  inv1 U996 ( .I(n893), .ZN(n66) );
  inv1 U997 ( .I(V116[10]), .ZN(n894) );
  or2 U998 ( .A1(n1529), .A2(n894), .Z(n895) );
  inv1 U999 ( .I(n895), .ZN(n63) );
  inv1 U1000 ( .I(V116[11]), .ZN(n896) );
  or2 U1001 ( .A1(n1529), .A2(n896), .Z(n897) );
  inv1 U1002 ( .I(n897), .ZN(n60) );
  inv1 U1003 ( .I(V116[12]), .ZN(n898) );
  or2 U1004 ( .A1(n1529), .A2(n898), .Z(n899) );
  inv1 U1005 ( .I(n899), .ZN(n57) );
  inv1 U1006 ( .I(V116[13]), .ZN(n900) );
  or2 U1007 ( .A1(n1529), .A2(n900), .Z(n901) );
  inv1 U1008 ( .I(n901), .ZN(n54) );
  inv1 U1009 ( .I(V116[14]), .ZN(n902) );
  or2 U1010 ( .A1(n1529), .A2(n902), .Z(n903) );
  inv1 U1011 ( .I(n903), .ZN(n51) );
  inv1 U1012 ( .I(V116[1]), .ZN(n904) );
  or2 U1013 ( .A1(n1529), .A2(n904), .Z(n905) );
  inv1 U1014 ( .I(n905), .ZN(n48) );
  inv1 U1015 ( .I(V116[2]), .ZN(n906) );
  or2 U1016 ( .A1(n1529), .A2(n906), .Z(n907) );
  inv1 U1017 ( .I(n907), .ZN(n45) );
  inv1 U1018 ( .I(V116[3]), .ZN(n908) );
  or2 U1019 ( .A1(n1529), .A2(n908), .Z(n909) );
  inv1 U1020 ( .I(n909), .ZN(n42) );
  inv1 U1021 ( .I(V116[4]), .ZN(n910) );
  or2 U1022 ( .A1(n1529), .A2(n910), .Z(n911) );
  inv1 U1023 ( .I(n911), .ZN(n39) );
  inv1 U1024 ( .I(V116[5]), .ZN(n912) );
  or2 U1025 ( .A1(n1529), .A2(n912), .Z(n913) );
  inv1 U1026 ( .I(n913), .ZN(n36) );
  inv1 U1027 ( .I(V116[6]), .ZN(n914) );
  or2 U1028 ( .A1(n1529), .A2(n914), .Z(n915) );
  inv1 U1029 ( .I(n915), .ZN(n33) );
  inv1 U1030 ( .I(V116[7]), .ZN(n916) );
  or2 U1031 ( .A1(n1529), .A2(n916), .Z(n917) );
  inv1 U1032 ( .I(n917), .ZN(n30) );
  inv1 U1033 ( .I(V116[8]), .ZN(n918) );
  or2 U1034 ( .A1(n1529), .A2(n918), .Z(n919) );
  inv1 U1035 ( .I(n919), .ZN(n27) );
  inv1 U1036 ( .I(V116[9]), .ZN(n920) );
  or2 U1037 ( .A1(n1529), .A2(n920), .Z(n921) );
  inv1 U1038 ( .I(n921), .ZN(n23) );
  inv1 U1039 ( .I(n930), .ZN(n929) );
  or2 U1040 ( .A1(n929), .A2(V133[8]), .Z(n924) );
  inv1 U1041 ( .I(n924), .ZN(n12) );
  and2 U1043 ( .A1(n1529), .A2(n1102), .Z(n926) );
  or2 U1044 ( .A1(n922), .A2(V119[0]), .Z(n923) );
  and2 U1045 ( .A1(n924), .A2(n923), .Z(n925) );
  and2 U1046 ( .A1(n926), .A2(n925), .Z(n10) );
  and2 U1047 ( .A1(n1738), .A2(n834), .Z(n927) );
  or2 U1048 ( .A1(n927), .A2(n7), .Z(n928) );
  and2 U1049 ( .A1(n929), .A2(n928), .Z(n1) );
  and2 U1050 ( .A1(V121[17]), .A2(n930), .Z(n2) );
  inv1 U1051 ( .I(n1101), .ZN(n1034) );
  inv1 U1052 ( .I(n981), .ZN(n931) );
  and2 U1053 ( .A1(n1739), .A2(n931), .Z(n932) );
  and2 U1054 ( .A1(n1034), .A2(n932), .Z(n933) );
  or2 U1055 ( .A1(n933), .A2(V133[10]), .Z(n934) );
  or2 U1056 ( .A1(n934), .A2(n752), .Z(n979) );
  or2 U1057 ( .A1(V133[6]), .A2(V133[5]), .Z(n954) );
  and2 U1058 ( .A1(n1739), .A2(n954), .Z(n936) );
  or2 U1059 ( .A1(n936), .A2(n853), .Z(n947) );
  inv1 U1060 ( .I(V133[3]), .ZN(n1072) );
  inv1 U1067 ( .I(V133[7]), .ZN(n955) );
  and2 U1068 ( .A1(n955), .A2(V133[5]), .Z(n942) );
  inv1 U1070 ( .I(n943), .ZN(n948) );
  and2 U1075 ( .A1(V15[0]), .A2(n1144), .Z(n953) );
  and2 U1076 ( .A1(n1102), .A2(n947), .Z(n951) );
  and2 U1081 ( .A1(V84[1]), .A2(n1141), .Z(n952) );
  or2 U1082 ( .A1(n953), .A2(n952), .Z(n962) );
  and2 U1083 ( .A1(n955), .A2(n954), .Z(n957) );
  or2 U1084 ( .A1(V133[1]), .A2(V133[2]), .Z(n956) );
  or2 U1085 ( .A1(n957), .A2(n956), .Z(n958) );
  inv1 U1086 ( .I(n958), .ZN(n959) );
  or2 U1089 ( .A1(n960), .A2(n1140), .Z(n961) );
  or2 U1090 ( .A1(n962), .A2(n961), .Z(n963) );
  and2 U1091 ( .A1(n979), .A2(n963), .Z(n972) );
  and2 U1092 ( .A1(V51[0]), .A2(n760), .Z(n965) );
  or2 U1093 ( .A1(n1739), .A2(n758), .Z(n984) );
  and2 U1094 ( .A1(n981), .A2(n984), .Z(n964) );
  and2 U1095 ( .A1(n965), .A2(n964), .Z(n970) );
  inv1 U1096 ( .I(n758), .ZN(n967) );
  and2 U1097 ( .A1(V50[0]), .A2(V133[8]), .Z(n966) );
  and2 U1098 ( .A1(n967), .A2(n966), .Z(n968) );
  or2 U1099 ( .A1(n968), .A2(n48), .Z(n969) );
  or2 U1100 ( .A1(n970), .A2(n969), .Z(n971) );
  or2 U1101 ( .A1(n972), .A2(n971), .Z(V136[0]) );
  or2 U1103 ( .A1(n973), .A2(n1140), .Z(n977) );
  and2 U1104 ( .A1(V84[2]), .A2(n1141), .Z(n975) );
  or2 U1106 ( .A1(n975), .A2(n974), .Z(n976) );
  or2 U1107 ( .A1(n977), .A2(n976), .Z(n978) );
  and2 U1108 ( .A1(n979), .A2(n978), .Z(n986) );
  and2 U1109 ( .A1(V52[0]), .A2(n760), .Z(n980) );
  and2 U1110 ( .A1(n981), .A2(n980), .Z(n982) );
  or2 U1111 ( .A1(n45), .A2(n982), .Z(n983) );
  and2 U1112 ( .A1(n984), .A2(n983), .Z(n985) );
  or2 U1113 ( .A1(n986), .A2(n985), .Z(V136[1]) );
  inv1 U1115 ( .I(n835), .ZN(n987) );
  or2 U1116 ( .A1(n1075), .A2(n987), .Z(n1063) );
  and2 U1117 ( .A1(V15[2]), .A2(n1144), .Z(n991) );
  and2 U1118 ( .A1(V47[3]), .A2(n855), .Z(n989) );
  and2 U1119 ( .A1(V84[3]), .A2(n1141), .Z(n988) );
  or2 U1120 ( .A1(n989), .A2(n988), .Z(n990) );
  or2 U1121 ( .A1(n991), .A2(n990), .Z(n992) );
  or2 U1123 ( .A1(n779), .A2(n42), .Z(n993) );
  or2 U1124 ( .A1(n994), .A2(n993), .Z(V142[0]) );
  and2 U1125 ( .A1(V15[3]), .A2(n1144), .Z(n998) );
  or2 U1128 ( .A1(n996), .A2(n995), .Z(n997) );
  or2 U1129 ( .A1(n998), .A2(n997), .Z(n999) );
  and2 U1130 ( .A1(n1063), .A2(n999), .Z(n1001) );
  or2 U1131 ( .A1(n779), .A2(n39), .Z(n1000) );
  and2 U1133 ( .A1(V15[4]), .A2(n1144), .Z(n1005) );
  or2 U1136 ( .A1(n1003), .A2(n1002), .Z(n1004) );
  or2 U1137 ( .A1(n1005), .A2(n1004), .Z(n1006) );
  and2 U1138 ( .A1(n1063), .A2(n1006), .Z(n1008) );
  or2 U1139 ( .A1(n779), .A2(n36), .Z(n1007) );
  or2 U1140 ( .A1(n1008), .A2(n1007), .Z(V142[2]) );
  and2 U1141 ( .A1(V15[5]), .A2(n1144), .Z(n1012) );
  and2 U1142 ( .A1(n855), .A2(V47[6]), .Z(n1010) );
  and2 U1143 ( .A1(V84[6]), .A2(n1141), .Z(n1009) );
  or2 U1144 ( .A1(n1010), .A2(n1009), .Z(n1011) );
  or2 U1145 ( .A1(n1012), .A2(n1011), .Z(n1013) );
  or2 U1147 ( .A1(n779), .A2(n33), .Z(n1014) );
  or2 U1148 ( .A1(n1015), .A2(n1014), .Z(V142[3]) );
  and2 U1149 ( .A1(V15[6]), .A2(n1144), .Z(n1020) );
  and2 U1150 ( .A1(V47[7]), .A2(n855), .Z(n1018) );
  and2 U1151 ( .A1(V84[7]), .A2(n1141), .Z(n1017) );
  or2 U1152 ( .A1(n1018), .A2(n1017), .Z(n1019) );
  or2 U1155 ( .A1(n779), .A2(n30), .Z(n1022) );
  or2 U1156 ( .A1(n1023), .A2(n1022), .Z(V142[4]) );
  and2 U1157 ( .A1(n1045), .A2(V47[0]), .Z(n1025) );
  and2 U1159 ( .A1(V84[8]), .A2(n1141), .Z(n1026) );
  or2 U1160 ( .A1(n1027), .A2(n1026), .Z(n1031) );
  and2 U1161 ( .A1(V15[7]), .A2(n1144), .Z(n1029) );
  and2 U1162 ( .A1(V47[8]), .A2(n856), .Z(n1028) );
  or2 U1163 ( .A1(n1029), .A2(n1028), .Z(n1030) );
  or2 U1164 ( .A1(n1031), .A2(n1030), .Z(n1032) );
  or2 U1166 ( .A1(n27), .A2(n1033), .Z(V142[5]) );
  or2 U1167 ( .A1(n1034), .A2(n1075), .Z(n1043) );
  or2 U1171 ( .A1(n1037), .A2(n1036), .Z(n1041) );
  and2 U1172 ( .A1(V15[8]), .A2(n1144), .Z(n1039) );
  and2 U1173 ( .A1(V47[9]), .A2(n856), .Z(n1038) );
  or2 U1174 ( .A1(n1039), .A2(n1038), .Z(n1040) );
  or2 U1175 ( .A1(n1041), .A2(n1040), .Z(n1042) );
  and2 U1176 ( .A1(n1043), .A2(n1042), .Z(n1044) );
  and2 U1179 ( .A1(n1045), .A2(V47[2]), .Z(n1046) );
  and2 U1181 ( .A1(V84[10]), .A2(n1141), .Z(n1047) );
  or2 U1182 ( .A1(n1048), .A2(n1047), .Z(n1052) );
  and2 U1183 ( .A1(V15[9]), .A2(n1144), .Z(n1050) );
  and2 U1184 ( .A1(V47[10]), .A2(n856), .Z(n1049) );
  or2 U1185 ( .A1(n1050), .A2(n1049), .Z(n1051) );
  and2 U1187 ( .A1(n1063), .A2(n1053), .Z(n1054) );
  or2 U1188 ( .A1(n63), .A2(n1054), .Z(V145[0]) );
  and2 U1189 ( .A1(n1045), .A2(V47[3]), .Z(n1055) );
  and2 U1191 ( .A1(V84[11]), .A2(n1141), .Z(n1056) );
  or2 U1192 ( .A1(n1057), .A2(n1056), .Z(n1061) );
  and2 U1193 ( .A1(V15[10]), .A2(n1144), .Z(n1059) );
  and2 U1194 ( .A1(V47[11]), .A2(n856), .Z(n1058) );
  or2 U1195 ( .A1(n1059), .A2(n1058), .Z(n1060) );
  or2 U1198 ( .A1(n60), .A2(n1064), .Z(V145[1]) );
  and2 U1199 ( .A1(n1045), .A2(V47[4]), .Z(n1065) );
  or2 U1200 ( .A1(n1140), .A2(n1065), .Z(n1067) );
  and2 U1201 ( .A1(V47[1]), .A2(n1141), .Z(n1066) );
  or2 U1202 ( .A1(n1067), .A2(n1066), .Z(n1071) );
  and2 U1203 ( .A1(V15[11]), .A2(n1144), .Z(n1069) );
  and2 U1204 ( .A1(V47[12]), .A2(n856), .Z(n1068) );
  or2 U1205 ( .A1(n1069), .A2(n1068), .Z(n1070) );
  or2 U1207 ( .A1(n836), .A2(n1072), .Z(n1073) );
  inv1 U1208 ( .I(n1073), .ZN(n1078) );
  inv1 U1210 ( .I(n1074), .ZN(n1076) );
  or2 U1213 ( .A1(n836), .A2(V133[1]), .Z(n1135) );
  inv1 U1214 ( .I(n1135), .ZN(n1079) );
  or2 U1215 ( .A1(n1090), .A2(n1079), .Z(n1080) );
  and2 U1217 ( .A1(V84[12]), .A2(n630), .Z(n1082) );
  and2 U1218 ( .A1(n834), .A2(n1082), .Z(n1084) );
  inv1 U1219 ( .I(V133[4]), .ZN(n1129) );
  and2 U1220 ( .A1(n1129), .A2(n1529), .Z(n1083) );
  and2 U1221 ( .A1(n1084), .A2(n1083), .Z(n1085) );
  or2 U1222 ( .A1(n57), .A2(n1085), .Z(n1086) );
  or2 U1223 ( .A1(n1087), .A2(n1086), .Z(V146[0]) );
  inv1 U1224 ( .I(n1088), .ZN(n1089) );
  or2 U1227 ( .A1(n1098), .A2(n832), .Z(n1091) );
  or2 U1228 ( .A1(n54), .A2(n859), .Z(n1096) );
  and2 U1230 ( .A1(n791), .A2(V47[5]), .Z(n1094) );
  and2 U1232 ( .A1(V47[2]), .A2(n865), .Z(n1093) );
  or2 U1233 ( .A1(n1094), .A2(n1093), .Z(n1095) );
  or2 U1234 ( .A1(n1096), .A2(n1095), .Z(n1107) );
  and2 U1236 ( .A1(V15[12]), .A2(n867), .Z(n1100) );
  and2 U1238 ( .A1(n868), .A2(V47[13]), .Z(n1099) );
  or2 U1239 ( .A1(n1100), .A2(n1099), .Z(n1105) );
  or2 U1240 ( .A1(n836), .A2(n631), .Z(n1103) );
  or2 U1241 ( .A1(n1103), .A2(n1102), .Z(n1309) );
  inv1 U1242 ( .I(n1309), .ZN(n1323) );
  and2 U1243 ( .A1(V84[13]), .A2(n1323), .Z(n1104) );
  or2 U1244 ( .A1(n1105), .A2(n1104), .Z(n1106) );
  or2 U1245 ( .A1(n1107), .A2(n1106), .Z(V149[0]) );
  or2 U1246 ( .A1(n51), .A2(n860), .Z(n1111) );
  and2 U1247 ( .A1(n791), .A2(V47[6]), .Z(n1109) );
  or2 U1249 ( .A1(n1109), .A2(n1108), .Z(n1110) );
  or2 U1250 ( .A1(n1111), .A2(n1110), .Z(n1117) );
  and2 U1251 ( .A1(V15[13]), .A2(n867), .Z(n1113) );
  and2 U1252 ( .A1(n868), .A2(V47[14]), .Z(n1112) );
  or2 U1253 ( .A1(n1113), .A2(n1112), .Z(n1115) );
  and2 U1254 ( .A1(V84[14]), .A2(n1323), .Z(n1114) );
  or2 U1255 ( .A1(n1115), .A2(n1114), .Z(n1116) );
  or2 U1256 ( .A1(n1117), .A2(n1116), .Z(V149[1]) );
  inv1 U1257 ( .I(V47[15]), .ZN(n1226) );
  inv1 U1259 ( .I(V84[15]), .ZN(n1711) );
  or2 U1260 ( .A1(n1309), .A2(n1711), .Z(n1118) );
  and2 U1261 ( .A1(n1119), .A2(n1118), .Z(n1121) );
  inv1 U1262 ( .I(V116[15]), .ZN(n1120) );
  or2 U1263 ( .A1(n1529), .A2(n1120), .Z(n1516) );
  and2 U1264 ( .A1(n1121), .A2(n1516), .Z(n1122) );
  inv1 U1265 ( .I(n1122), .ZN(n1128) );
  and2 U1266 ( .A1(V15[14]), .A2(n867), .Z(n1124) );
  and2 U1267 ( .A1(V47[4]), .A2(n865), .Z(n1123) );
  or2 U1268 ( .A1(n1124), .A2(n1123), .Z(n1126) );
  or2 U1269 ( .A1(n787), .A2(n859), .Z(n1125) );
  or2 U1270 ( .A1(n1126), .A2(n1125), .Z(n1127) );
  or2 U1271 ( .A1(n1128), .A2(n1127), .Z(V149[2]) );
  and2 U1272 ( .A1(V84[16]), .A2(n630), .Z(n1131) );
  and2 U1273 ( .A1(n1129), .A2(n834), .Z(n1130) );
  and2 U1274 ( .A1(n1131), .A2(n1130), .Z(n1132) );
  or2 U1275 ( .A1(n872), .A2(n1132), .Z(n1134) );
  or2 U1276 ( .A1(V116[16]), .A2(n1529), .Z(n1133) );
  and2 U1277 ( .A1(n1134), .A2(n1133), .Z(n1152) );
  or2 U1278 ( .A1(V133[2]), .A2(n1135), .Z(n1137) );
  and2 U1279 ( .A1(n1137), .A2(n1098), .Z(n1138) );
  inv1 U1280 ( .I(n1138), .ZN(n1150) );
  or2 U1282 ( .A1(n1140), .A2(n1139), .Z(n1143) );
  or2 U1284 ( .A1(n1143), .A2(n1142), .Z(n1148) );
  and2 U1285 ( .A1(V47[1]), .A2(n1144), .Z(n1146) );
  and2 U1286 ( .A1(V47[16]), .A2(n856), .Z(n1145) );
  or2 U1287 ( .A1(n1146), .A2(n1145), .Z(n1147) );
  or2 U1288 ( .A1(n1148), .A2(n1147), .Z(n1149) );
  and2 U1289 ( .A1(n1150), .A2(n1149), .Z(n1151) );
  inv1 U1291 ( .I(V47[17]), .ZN(n1352) );
  inv1 U1293 ( .I(V84[17]), .ZN(n1644) );
  or2 U1294 ( .A1(n1309), .A2(n1644), .Z(n1153) );
  and2 U1295 ( .A1(n1154), .A2(n1153), .Z(n1156) );
  inv1 U1296 ( .I(V116[17]), .ZN(n1155) );
  or2 U1297 ( .A1(n1529), .A2(n1155), .Z(n1541) );
  and2 U1298 ( .A1(n1156), .A2(n1541), .Z(n1157) );
  inv1 U1299 ( .I(n1157), .ZN(n1163) );
  and2 U1300 ( .A1(V47[2]), .A2(n867), .Z(n1159) );
  and2 U1301 ( .A1(V47[6]), .A2(n865), .Z(n1158) );
  or2 U1302 ( .A1(n1159), .A2(n1158), .Z(n1161) );
  or2 U1303 ( .A1(n789), .A2(n859), .Z(n1160) );
  or2 U1304 ( .A1(n1161), .A2(n1160), .Z(n1162) );
  or2 U1305 ( .A1(n1163), .A2(n1162), .Z(V165[0]) );
  inv1 U1306 ( .I(V47[18]), .ZN(n1368) );
  or2 U1307 ( .A1(n870), .A2(n1368), .Z(n1165) );
  inv1 U1308 ( .I(V84[18]), .ZN(n1659) );
  or2 U1309 ( .A1(n1309), .A2(n1659), .Z(n1164) );
  and2 U1310 ( .A1(n1165), .A2(n1164), .Z(n1167) );
  inv1 U1311 ( .I(V116[18]), .ZN(n1166) );
  or2 U1312 ( .A1(n1529), .A2(n1166), .Z(n1554) );
  and2 U1313 ( .A1(n1167), .A2(n1554), .Z(n1168) );
  inv1 U1314 ( .I(n1168), .ZN(n1174) );
  and2 U1315 ( .A1(V47[3]), .A2(n867), .Z(n1170) );
  and2 U1316 ( .A1(V47[7]), .A2(n866), .Z(n1169) );
  or2 U1317 ( .A1(n1170), .A2(n1169), .Z(n1172) );
  or2 U1318 ( .A1(n790), .A2(n860), .Z(n1171) );
  or2 U1319 ( .A1(n1172), .A2(n1171), .Z(n1173) );
  or2 U1320 ( .A1(n1174), .A2(n1173), .Z(V165[1]) );
  inv1 U1321 ( .I(V47[19]), .ZN(n1379) );
  or2 U1322 ( .A1(n871), .A2(n1379), .Z(n1176) );
  inv1 U1323 ( .I(V84[19]), .ZN(n1674) );
  or2 U1324 ( .A1(n1309), .A2(n1674), .Z(n1175) );
  and2 U1325 ( .A1(n1176), .A2(n1175), .Z(n1178) );
  inv1 U1326 ( .I(V116[19]), .ZN(n1177) );
  or2 U1327 ( .A1(n1529), .A2(n1177), .Z(n1566) );
  and2 U1328 ( .A1(n1178), .A2(n1566), .Z(n1179) );
  inv1 U1329 ( .I(n1179), .ZN(n1185) );
  and2 U1330 ( .A1(V47[4]), .A2(n867), .Z(n1181) );
  and2 U1331 ( .A1(V47[8]), .A2(n866), .Z(n1180) );
  or2 U1332 ( .A1(n1181), .A2(n1180), .Z(n1183) );
  or2 U1333 ( .A1(n792), .A2(n860), .Z(n1182) );
  or2 U1334 ( .A1(n1183), .A2(n1182), .Z(n1184) );
  or2 U1335 ( .A1(n1185), .A2(n1184), .Z(V165[2]) );
  inv1 U1336 ( .I(V47[20]), .ZN(n1390) );
  inv1 U1338 ( .I(V84[20]), .ZN(n1689) );
  or2 U1339 ( .A1(n1309), .A2(n1689), .Z(n1186) );
  and2 U1340 ( .A1(n1187), .A2(n1186), .Z(n1189) );
  inv1 U1341 ( .I(V116[20]), .ZN(n1188) );
  or2 U1342 ( .A1(n1529), .A2(n1188), .Z(n1577) );
  and2 U1343 ( .A1(n1189), .A2(n1577), .Z(n1190) );
  inv1 U1344 ( .I(n1190), .ZN(n1196) );
  and2 U1345 ( .A1(V47[5]), .A2(n867), .Z(n1192) );
  and2 U1346 ( .A1(V47[9]), .A2(n865), .Z(n1191) );
  or2 U1347 ( .A1(n1192), .A2(n1191), .Z(n1194) );
  or2 U1348 ( .A1(n794), .A2(n859), .Z(n1193) );
  or2 U1349 ( .A1(n1194), .A2(n1193), .Z(n1195) );
  or2 U1350 ( .A1(n1196), .A2(n1195), .Z(V165[3]) );
  inv1 U1351 ( .I(V47[21]), .ZN(n1401) );
  or2 U1352 ( .A1(n870), .A2(n1401), .Z(n1198) );
  inv1 U1353 ( .I(V84[21]), .ZN(n1704) );
  or2 U1354 ( .A1(n1309), .A2(n1704), .Z(n1197) );
  and2 U1355 ( .A1(n1198), .A2(n1197), .Z(n1200) );
  inv1 U1356 ( .I(V116[21]), .ZN(n1199) );
  or2 U1357 ( .A1(n1529), .A2(n1199), .Z(n1590) );
  and2 U1358 ( .A1(n1200), .A2(n1590), .Z(n1201) );
  inv1 U1359 ( .I(n1201), .ZN(n1207) );
  and2 U1360 ( .A1(V47[6]), .A2(n867), .Z(n1203) );
  and2 U1361 ( .A1(V47[10]), .A2(n866), .Z(n1202) );
  or2 U1362 ( .A1(n1203), .A2(n1202), .Z(n1205) );
  or2 U1363 ( .A1(n795), .A2(n860), .Z(n1204) );
  or2 U1364 ( .A1(n1205), .A2(n1204), .Z(n1206) );
  or2 U1365 ( .A1(n1207), .A2(n1206), .Z(V165[4]) );
  inv1 U1366 ( .I(V47[22]), .ZN(n1410) );
  or2 U1367 ( .A1(n871), .A2(n1410), .Z(n1209) );
  inv1 U1368 ( .I(V84[22]), .ZN(n1719) );
  or2 U1369 ( .A1(n1309), .A2(n1719), .Z(n1208) );
  and2 U1370 ( .A1(n1209), .A2(n1208), .Z(n1211) );
  inv1 U1371 ( .I(V116[22]), .ZN(n1210) );
  or2 U1372 ( .A1(n1529), .A2(n1210), .Z(n1601) );
  and2 U1373 ( .A1(n1211), .A2(n1601), .Z(n1212) );
  inv1 U1374 ( .I(n1212), .ZN(n1218) );
  and2 U1375 ( .A1(V47[7]), .A2(n867), .Z(n1214) );
  and2 U1376 ( .A1(V47[11]), .A2(n865), .Z(n1213) );
  or2 U1377 ( .A1(n1214), .A2(n1213), .Z(n1216) );
  or2 U1378 ( .A1(n796), .A2(n860), .Z(n1215) );
  or2 U1379 ( .A1(n1216), .A2(n1215), .Z(n1217) );
  or2 U1380 ( .A1(n1218), .A2(n1217), .Z(V165[5]) );
  inv1 U1381 ( .I(V47[23]), .ZN(n1421) );
  or2 U1382 ( .A1(n870), .A2(n1421), .Z(n1220) );
  inv1 U1383 ( .I(V84[23]), .ZN(n1608) );
  or2 U1384 ( .A1(n1309), .A2(n1608), .Z(n1219) );
  and2 U1385 ( .A1(n1220), .A2(n1219), .Z(n1222) );
  inv1 U1386 ( .I(V116[23]), .ZN(n1221) );
  or2 U1387 ( .A1(n1529), .A2(n1221), .Z(n1612) );
  and2 U1388 ( .A1(n1222), .A2(n1612), .Z(n1223) );
  inv1 U1389 ( .I(n1223), .ZN(n1232) );
  and2 U1390 ( .A1(V47[8]), .A2(n867), .Z(n1225) );
  and2 U1391 ( .A1(V47[12]), .A2(n865), .Z(n1224) );
  or2 U1392 ( .A1(n1225), .A2(n1224), .Z(n1230) );
  or2 U1393 ( .A1(n863), .A2(n1226), .Z(n1227) );
  inv1 U1394 ( .I(n1227), .ZN(n1228) );
  or2 U1395 ( .A1(n1228), .A2(n859), .Z(n1229) );
  or2 U1396 ( .A1(n1230), .A2(n1229), .Z(n1231) );
  or2 U1397 ( .A1(n1232), .A2(n1231), .Z(V165[6]) );
  inv1 U1398 ( .I(V47[24]), .ZN(n1432) );
  or2 U1399 ( .A1(n871), .A2(n1432), .Z(n1234) );
  inv1 U1400 ( .I(V84[24]), .ZN(n1622) );
  or2 U1401 ( .A1(n1309), .A2(n1622), .Z(n1233) );
  and2 U1402 ( .A1(n1234), .A2(n1233), .Z(n1236) );
  inv1 U1403 ( .I(V116[24]), .ZN(n1235) );
  or2 U1404 ( .A1(n1529), .A2(n1235), .Z(n1626) );
  and2 U1405 ( .A1(n1236), .A2(n1626), .Z(n1237) );
  inv1 U1406 ( .I(n1237), .ZN(n1243) );
  and2 U1407 ( .A1(V47[9]), .A2(n867), .Z(n1239) );
  and2 U1408 ( .A1(V47[13]), .A2(n866), .Z(n1238) );
  or2 U1409 ( .A1(n1239), .A2(n1238), .Z(n1241) );
  or2 U1410 ( .A1(n798), .A2(n860), .Z(n1240) );
  or2 U1411 ( .A1(n1241), .A2(n1240), .Z(n1242) );
  or2 U1412 ( .A1(n1243), .A2(n1242), .Z(V165[7]) );
  inv1 U1413 ( .I(V47[25]), .ZN(n1441) );
  or2 U1414 ( .A1(n871), .A2(n1441), .Z(n1245) );
  inv1 U1415 ( .I(V84[25]), .ZN(n1637) );
  or2 U1416 ( .A1(n1309), .A2(n1637), .Z(n1244) );
  and2 U1417 ( .A1(n1245), .A2(n1244), .Z(n1247) );
  inv1 U1418 ( .I(V116[25]), .ZN(n1246) );
  or2 U1419 ( .A1(n1529), .A2(n1246), .Z(n1641) );
  and2 U1420 ( .A1(n1247), .A2(n1641), .Z(n1248) );
  inv1 U1421 ( .I(n1248), .ZN(n1256) );
  and2 U1422 ( .A1(V47[10]), .A2(n867), .Z(n1250) );
  and2 U1423 ( .A1(V47[14]), .A2(n865), .Z(n1249) );
  or2 U1424 ( .A1(n1250), .A2(n1249), .Z(n1254) );
  or2 U1425 ( .A1(n863), .A2(n1352), .Z(n1251) );
  inv1 U1426 ( .I(n1251), .ZN(n1252) );
  or2 U1427 ( .A1(n1252), .A2(n859), .Z(n1253) );
  or2 U1428 ( .A1(n1254), .A2(n1253), .Z(n1255) );
  or2 U1429 ( .A1(n1256), .A2(n1255), .Z(V165[8]) );
  inv1 U1430 ( .I(V47[26]), .ZN(n1452) );
  inv1 U1432 ( .I(V84[26]), .ZN(n1652) );
  or2 U1433 ( .A1(n1309), .A2(n1652), .Z(n1257) );
  and2 U1434 ( .A1(n1258), .A2(n1257), .Z(n1260) );
  inv1 U1435 ( .I(V116[26]), .ZN(n1259) );
  or2 U1436 ( .A1(n1529), .A2(n1259), .Z(n1656) );
  and2 U1437 ( .A1(n1260), .A2(n1656), .Z(n1261) );
  inv1 U1438 ( .I(n1261), .ZN(n1269) );
  and2 U1439 ( .A1(V47[11]), .A2(n867), .Z(n1263) );
  and2 U1440 ( .A1(V47[15]), .A2(n865), .Z(n1262) );
  or2 U1441 ( .A1(n1263), .A2(n1262), .Z(n1267) );
  or2 U1442 ( .A1(n864), .A2(n1368), .Z(n1264) );
  inv1 U1443 ( .I(n1264), .ZN(n1265) );
  or2 U1444 ( .A1(n1265), .A2(n859), .Z(n1266) );
  or2 U1445 ( .A1(n1267), .A2(n1266), .Z(n1268) );
  or2 U1446 ( .A1(n1269), .A2(n1268), .Z(V165[9]) );
  inv1 U1447 ( .I(V47[27]), .ZN(n1461) );
  or2 U1448 ( .A1(n870), .A2(n1461), .Z(n1271) );
  inv1 U1449 ( .I(V84[27]), .ZN(n1667) );
  or2 U1450 ( .A1(n1309), .A2(n1667), .Z(n1270) );
  and2 U1451 ( .A1(n1271), .A2(n1270), .Z(n1273) );
  inv1 U1452 ( .I(V116[27]), .ZN(n1272) );
  or2 U1453 ( .A1(n1529), .A2(n1272), .Z(n1671) );
  and2 U1454 ( .A1(n1273), .A2(n1671), .Z(n1274) );
  inv1 U1455 ( .I(n1274), .ZN(n1282) );
  and2 U1456 ( .A1(V47[12]), .A2(n867), .Z(n1276) );
  and2 U1457 ( .A1(V47[16]), .A2(n866), .Z(n1275) );
  or2 U1458 ( .A1(n1276), .A2(n1275), .Z(n1280) );
  or2 U1459 ( .A1(n864), .A2(n1379), .Z(n1277) );
  inv1 U1460 ( .I(n1277), .ZN(n1278) );
  or2 U1461 ( .A1(n1278), .A2(n860), .Z(n1279) );
  or2 U1462 ( .A1(n1280), .A2(n1279), .Z(n1281) );
  or2 U1463 ( .A1(n1282), .A2(n1281), .Z(V165[10]) );
  inv1 U1464 ( .I(V47[28]), .ZN(n1472) );
  or2 U1465 ( .A1(n870), .A2(n1472), .Z(n1284) );
  inv1 U1466 ( .I(V84[28]), .ZN(n1682) );
  or2 U1467 ( .A1(n1309), .A2(n1682), .Z(n1283) );
  and2 U1468 ( .A1(n1284), .A2(n1283), .Z(n1286) );
  inv1 U1469 ( .I(V116[28]), .ZN(n1285) );
  or2 U1470 ( .A1(n1529), .A2(n1285), .Z(n1686) );
  and2 U1471 ( .A1(n1286), .A2(n1686), .Z(n1287) );
  inv1 U1472 ( .I(n1287), .ZN(n1295) );
  and2 U1473 ( .A1(V47[13]), .A2(n867), .Z(n1289) );
  and2 U1474 ( .A1(V47[17]), .A2(n866), .Z(n1288) );
  or2 U1475 ( .A1(n1289), .A2(n1288), .Z(n1293) );
  or2 U1476 ( .A1(n864), .A2(n1390), .Z(n1290) );
  inv1 U1477 ( .I(n1290), .ZN(n1291) );
  or2 U1478 ( .A1(n1291), .A2(n860), .Z(n1292) );
  or2 U1479 ( .A1(n1293), .A2(n1292), .Z(n1294) );
  or2 U1480 ( .A1(n1295), .A2(n1294), .Z(V165[11]) );
  inv1 U1481 ( .I(V47[29]), .ZN(n1481) );
  or2 U1482 ( .A1(n871), .A2(n1481), .Z(n1297) );
  inv1 U1483 ( .I(V84[29]), .ZN(n1697) );
  or2 U1484 ( .A1(n1309), .A2(n1697), .Z(n1296) );
  and2 U1485 ( .A1(n1297), .A2(n1296), .Z(n1299) );
  inv1 U1486 ( .I(V116[29]), .ZN(n1298) );
  or2 U1487 ( .A1(n1529), .A2(n1298), .Z(n1701) );
  and2 U1488 ( .A1(n1299), .A2(n1701), .Z(n1300) );
  inv1 U1489 ( .I(n1300), .ZN(n1308) );
  and2 U1490 ( .A1(V47[14]), .A2(n867), .Z(n1302) );
  and2 U1491 ( .A1(V47[18]), .A2(n865), .Z(n1301) );
  or2 U1492 ( .A1(n1302), .A2(n1301), .Z(n1306) );
  or2 U1493 ( .A1(n864), .A2(n1401), .Z(n1303) );
  inv1 U1494 ( .I(n1303), .ZN(n1304) );
  or2 U1495 ( .A1(n1304), .A2(n859), .Z(n1305) );
  or2 U1496 ( .A1(n1306), .A2(n1305), .Z(n1307) );
  or2 U1497 ( .A1(n1308), .A2(n1307), .Z(V165[12]) );
  inv1 U1498 ( .I(V47[30]), .ZN(n1492) );
  inv1 U1500 ( .I(V84[30]), .ZN(n1712) );
  or2 U1501 ( .A1(n1309), .A2(n1712), .Z(n1310) );
  and2 U1502 ( .A1(n1311), .A2(n1310), .Z(n1313) );
  inv1 U1503 ( .I(V116[30]), .ZN(n1312) );
  or2 U1504 ( .A1(n1529), .A2(n1312), .Z(n1716) );
  and2 U1505 ( .A1(n1313), .A2(n1716), .Z(n1314) );
  and2 U1507 ( .A1(V47[15]), .A2(n867), .Z(n1316) );
  and2 U1508 ( .A1(V47[19]), .A2(n866), .Z(n1315) );
  or2 U1509 ( .A1(n1316), .A2(n1315), .Z(n1320) );
  or2 U1510 ( .A1(n863), .A2(n1410), .Z(n1317) );
  inv1 U1511 ( .I(n1317), .ZN(n1318) );
  or2 U1512 ( .A1(n1318), .A2(n860), .Z(n1319) );
  or2 U1513 ( .A1(n1320), .A2(n1319), .Z(n1321) );
  or2 U1514 ( .A1(n1322), .A2(n1321), .Z(V165[13]) );
  and2 U1515 ( .A1(V84[31]), .A2(n1323), .Z(n1326) );
  inv1 U1516 ( .I(V116[31]), .ZN(n1324) );
  or2 U1517 ( .A1(n1529), .A2(n1324), .Z(n1325) );
  inv1 U1518 ( .I(n1325), .ZN(n1734) );
  or2 U1519 ( .A1(n1326), .A2(n1734), .Z(n1327) );
  or2 U1520 ( .A1(n1327), .A2(n859), .Z(n1339) );
  inv1 U1521 ( .I(V47[31]), .ZN(n1503) );
  or2 U1522 ( .A1(n871), .A2(n1503), .Z(n1329) );
  inv1 U1523 ( .I(n1329), .ZN(n1331) );
  and2 U1526 ( .A1(V47[20]), .A2(n866), .Z(n1335) );
  or2 U1527 ( .A1(n862), .A2(n1421), .Z(n1333) );
  inv1 U1528 ( .I(n1333), .ZN(n1334) );
  or2 U1529 ( .A1(n1335), .A2(n1334), .Z(n1336) );
  or2 U1530 ( .A1(n1337), .A2(n1336), .Z(n1338) );
  or2 U1531 ( .A1(n1339), .A2(n1338), .Z(V165[14]) );
  or2 U1534 ( .A1(n1342), .A2(V133[0]), .Z(n1343) );
  inv1 U1537 ( .I(n382), .ZN(n1348) );
  inv1 U1538 ( .I(n395), .ZN(n1347) );
  inv1 U1544 ( .I(V84[0]), .ZN(n1512) );
  or2 U1545 ( .A1(n1743), .A2(n1512), .Z(n1353) );
  and2 U1546 ( .A1(n1354), .A2(n1353), .Z(n1355) );
  inv1 U1547 ( .I(n1355), .ZN(n1356) );
  or2 U1548 ( .A1(n1356), .A2(n66), .Z(n1367) );
  and2 U1550 ( .A1(V47[21]), .A2(n876), .Z(n1365) );
  or2 U1552 ( .A1(n1753), .A2(n1432), .Z(n1359) );
  inv1 U1553 ( .I(n1359), .ZN(n1363) );
  or2 U1555 ( .A1(n1363), .A2(n883), .Z(n1364) );
  or2 U1556 ( .A1(n1364), .A2(n1365), .Z(n1366) );
  or2 U1557 ( .A1(n1367), .A2(n1366), .Z(V197[0]) );
  inv1 U1559 ( .I(V84[1]), .ZN(n1525) );
  or2 U1560 ( .A1(n1745), .A2(n1525), .Z(n1369) );
  and2 U1561 ( .A1(n1370), .A2(n1369), .Z(n1371) );
  inv1 U1562 ( .I(n1371), .ZN(n1372) );
  or2 U1563 ( .A1(n1372), .A2(n48), .Z(n1378) );
  and2 U1564 ( .A1(V47[22]), .A2(n876), .Z(n1376) );
  or2 U1565 ( .A1(n1753), .A2(n1441), .Z(n1373) );
  inv1 U1566 ( .I(n1373), .ZN(n1374) );
  or2 U1567 ( .A1(n1374), .A2(n882), .Z(n1375) );
  or2 U1568 ( .A1(n1375), .A2(n1376), .Z(n1377) );
  or2 U1569 ( .A1(n1378), .A2(n1377), .Z(V197[1]) );
  inv1 U1571 ( .I(V84[2]), .ZN(n1537) );
  or2 U1572 ( .A1(n1746), .A2(n1537), .Z(n1380) );
  and2 U1573 ( .A1(n1381), .A2(n1380), .Z(n1382) );
  inv1 U1574 ( .I(n1382), .ZN(n1383) );
  or2 U1575 ( .A1(n1383), .A2(n45), .Z(n1389) );
  and2 U1576 ( .A1(V47[23]), .A2(n1741), .Z(n1387) );
  or2 U1577 ( .A1(n1752), .A2(n1452), .Z(n1384) );
  inv1 U1578 ( .I(n1384), .ZN(n1385) );
  or2 U1579 ( .A1(n1385), .A2(n881), .Z(n1386) );
  or2 U1580 ( .A1(n1386), .A2(n1387), .Z(n1388) );
  or2 U1581 ( .A1(n1389), .A2(n1388), .Z(V197[2]) );
  or2 U1582 ( .A1(n844), .A2(n1390), .Z(n1392) );
  inv1 U1583 ( .I(V84[3]), .ZN(n1550) );
  or2 U1584 ( .A1(n1747), .A2(n1550), .Z(n1391) );
  and2 U1585 ( .A1(n1392), .A2(n1391), .Z(n1393) );
  or2 U1587 ( .A1(n1394), .A2(n42), .Z(n1400) );
  and2 U1588 ( .A1(V47[24]), .A2(n876), .Z(n1398) );
  or2 U1589 ( .A1(n1748), .A2(n1461), .Z(n1395) );
  inv1 U1590 ( .I(n1395), .ZN(n1396) );
  or2 U1591 ( .A1(n1396), .A2(n883), .Z(n1397) );
  or2 U1592 ( .A1(n1397), .A2(n1398), .Z(n1399) );
  or2 U1593 ( .A1(n1400), .A2(n1399), .Z(V197[3]) );
  inv1 U1595 ( .I(V84[4]), .ZN(n1562) );
  or2 U1596 ( .A1(n1744), .A2(n1562), .Z(n1402) );
  or2 U1597 ( .A1(n826), .A2(n39), .Z(n1409) );
  and2 U1598 ( .A1(V47[25]), .A2(n876), .Z(n1407) );
  or2 U1599 ( .A1(n1751), .A2(n1472), .Z(n1404) );
  inv1 U1600 ( .I(n1404), .ZN(n1405) );
  or2 U1601 ( .A1(n1405), .A2(n882), .Z(n1406) );
  or2 U1602 ( .A1(n1406), .A2(n1407), .Z(n1408) );
  or2 U1603 ( .A1(n1409), .A2(n1408), .Z(V197[4]) );
  inv1 U1605 ( .I(V84[5]), .ZN(n1573) );
  or2 U1606 ( .A1(n1744), .A2(n1573), .Z(n1411) );
  and2 U1607 ( .A1(n1412), .A2(n1411), .Z(n1413) );
  inv1 U1608 ( .I(n1413), .ZN(n1414) );
  or2 U1609 ( .A1(n1414), .A2(n36), .Z(n1420) );
  and2 U1610 ( .A1(V47[26]), .A2(n876), .Z(n1418) );
  or2 U1611 ( .A1(n1752), .A2(n1481), .Z(n1415) );
  inv1 U1612 ( .I(n1415), .ZN(n1416) );
  or2 U1613 ( .A1(n1416), .A2(n883), .Z(n1417) );
  or2 U1614 ( .A1(n1417), .A2(n1418), .Z(n1419) );
  or2 U1615 ( .A1(n1420), .A2(n1419), .Z(V197[5]) );
  inv1 U1617 ( .I(V84[6]), .ZN(n1586) );
  or2 U1618 ( .A1(n1745), .A2(n1586), .Z(n1422) );
  inv1 U1620 ( .I(n1424), .ZN(n1425) );
  or2 U1621 ( .A1(n1425), .A2(n33), .Z(n1431) );
  and2 U1622 ( .A1(V47[27]), .A2(n876), .Z(n1429) );
  or2 U1623 ( .A1(n1749), .A2(n1492), .Z(n1426) );
  inv1 U1624 ( .I(n1426), .ZN(n1427) );
  or2 U1625 ( .A1(n1427), .A2(n881), .Z(n1428) );
  or2 U1626 ( .A1(n1428), .A2(n1429), .Z(n1430) );
  or2 U1627 ( .A1(n1431), .A2(n1430), .Z(V197[6]) );
  or2 U1628 ( .A1(n844), .A2(n1432), .Z(n1434) );
  inv1 U1629 ( .I(V84[7]), .ZN(n1598) );
  or2 U1630 ( .A1(n1746), .A2(n1598), .Z(n1433) );
  or2 U1631 ( .A1(n827), .A2(n30), .Z(n1440) );
  and2 U1632 ( .A1(V47[28]), .A2(n875), .Z(n1438) );
  or2 U1633 ( .A1(n1753), .A2(n1503), .Z(n1435) );
  inv1 U1634 ( .I(n1435), .ZN(n1436) );
  or2 U1635 ( .A1(n1436), .A2(n883), .Z(n1437) );
  or2 U1636 ( .A1(n1437), .A2(n1438), .Z(n1439) );
  or2 U1637 ( .A1(n1440), .A2(n1439), .Z(V197[7]) );
  or2 U1638 ( .A1(n805), .A2(n1441), .Z(n1443) );
  inv1 U1639 ( .I(V84[8]), .ZN(n1607) );
  or2 U1640 ( .A1(n1744), .A2(n1607), .Z(n1442) );
  or2 U1643 ( .A1(n1445), .A2(n27), .Z(n1451) );
  and2 U1644 ( .A1(V47[29]), .A2(n875), .Z(n1449) );
  or2 U1645 ( .A1(n1751), .A2(n1512), .Z(n1446) );
  inv1 U1646 ( .I(n1446), .ZN(n1447) );
  or2 U1647 ( .A1(n1447), .A2(n882), .Z(n1448) );
  or2 U1648 ( .A1(n1448), .A2(n1449), .Z(n1450) );
  or2 U1649 ( .A1(n1451), .A2(n1450), .Z(V197[8]) );
  inv1 U1651 ( .I(V84[9]), .ZN(n1621) );
  or2 U1652 ( .A1(n1743), .A2(n1621), .Z(n1453) );
  or2 U1655 ( .A1(n1456), .A2(n23), .Z(n1460) );
  and2 U1656 ( .A1(V47[30]), .A2(n876), .Z(n1458) );
  or2 U1657 ( .A1(n810), .A2(n881), .Z(n1457) );
  or2 U1658 ( .A1(n1457), .A2(n1458), .Z(n1459) );
  or2 U1659 ( .A1(n1460), .A2(n1459), .Z(V197[9]) );
  inv1 U1661 ( .I(V84[10]), .ZN(n1636) );
  or2 U1662 ( .A1(n1747), .A2(n1636), .Z(n1462) );
  inv1 U1664 ( .I(n1464), .ZN(n1465) );
  or2 U1665 ( .A1(n1465), .A2(n63), .Z(n1471) );
  and2 U1666 ( .A1(V47[31]), .A2(n875), .Z(n1469) );
  or2 U1667 ( .A1(n1749), .A2(n1537), .Z(n1466) );
  inv1 U1668 ( .I(n1466), .ZN(n1467) );
  or2 U1669 ( .A1(n1467), .A2(n882), .Z(n1468) );
  or2 U1670 ( .A1(n1469), .A2(n1468), .Z(n1470) );
  or2 U1671 ( .A1(n1471), .A2(n1470), .Z(V197[10]) );
  inv1 U1673 ( .I(V84[11]), .ZN(n1651) );
  or2 U1674 ( .A1(n1745), .A2(n1651), .Z(n1473) );
  or2 U1675 ( .A1(n846), .A2(n60), .Z(n1480) );
  and2 U1676 ( .A1(V84[0]), .A2(n875), .Z(n1478) );
  or2 U1677 ( .A1(n1749), .A2(n1550), .Z(n1475) );
  inv1 U1678 ( .I(n1475), .ZN(n1476) );
  or2 U1679 ( .A1(n1476), .A2(n881), .Z(n1477) );
  or2 U1680 ( .A1(n1477), .A2(n1478), .Z(n1479) );
  or2 U1681 ( .A1(n1480), .A2(n1479), .Z(V197[11]) );
  inv1 U1683 ( .I(V84[12]), .ZN(n1666) );
  or2 U1684 ( .A1(n1746), .A2(n1666), .Z(n1482) );
  and2 U1685 ( .A1(n1483), .A2(n1482), .Z(n1484) );
  inv1 U1686 ( .I(n1484), .ZN(n1485) );
  or2 U1687 ( .A1(n1485), .A2(n57), .Z(n1491) );
  and2 U1688 ( .A1(V84[1]), .A2(n1741), .Z(n1489) );
  or2 U1689 ( .A1(n1749), .A2(n1562), .Z(n1486) );
  inv1 U1690 ( .I(n1486), .ZN(n1487) );
  or2 U1691 ( .A1(n1487), .A2(n883), .Z(n1488) );
  or2 U1692 ( .A1(n1488), .A2(n1489), .Z(n1490) );
  or2 U1693 ( .A1(n1491), .A2(n1490), .Z(V197[12]) );
  inv1 U1695 ( .I(V84[13]), .ZN(n1681) );
  or2 U1696 ( .A1(n1743), .A2(n1681), .Z(n1493) );
  and2 U1697 ( .A1(n1494), .A2(n1493), .Z(n1495) );
  inv1 U1698 ( .I(n1495), .ZN(n1496) );
  or2 U1699 ( .A1(n1496), .A2(n54), .Z(n1502) );
  and2 U1700 ( .A1(V84[2]), .A2(n876), .Z(n1500) );
  or2 U1701 ( .A1(n1750), .A2(n1573), .Z(n1497) );
  inv1 U1702 ( .I(n1497), .ZN(n1498) );
  or2 U1703 ( .A1(n1498), .A2(n883), .Z(n1499) );
  or2 U1704 ( .A1(n1499), .A2(n1500), .Z(n1501) );
  or2 U1705 ( .A1(n1502), .A2(n1501), .Z(V197[13]) );
  inv1 U1707 ( .I(V84[14]), .ZN(n1696) );
  or2 U1708 ( .A1(n1744), .A2(n1696), .Z(n1504) );
  or2 U1709 ( .A1(n820), .A2(n51), .Z(n1511) );
  and2 U1710 ( .A1(V84[3]), .A2(n876), .Z(n1509) );
  or2 U1711 ( .A1(n1752), .A2(n1586), .Z(n1506) );
  inv1 U1712 ( .I(n1506), .ZN(n1507) );
  or2 U1713 ( .A1(n1507), .A2(n881), .Z(n1508) );
  or2 U1714 ( .A1(n1508), .A2(n1509), .Z(n1510) );
  or2 U1715 ( .A1(n1511), .A2(n1510), .Z(V197[14]) );
  or2 U1717 ( .A1(n1744), .A2(n1711), .Z(n1513) );
  and2 U1718 ( .A1(n1514), .A2(n1513), .Z(n1515) );
  inv1 U1719 ( .I(n1515), .ZN(n1518) );
  inv1 U1720 ( .I(n1516), .ZN(n1517) );
  or2 U1721 ( .A1(n1518), .A2(n1517), .Z(n1524) );
  and2 U1722 ( .A1(V84[4]), .A2(n875), .Z(n1522) );
  or2 U1723 ( .A1(n1751), .A2(n1598), .Z(n1519) );
  inv1 U1724 ( .I(n1519), .ZN(n1520) );
  or2 U1725 ( .A1(n1520), .A2(n883), .Z(n1521) );
  or2 U1726 ( .A1(n1521), .A2(n1522), .Z(n1523) );
  or2 U1727 ( .A1(n1524), .A2(n1523), .Z(V197[15]) );
  inv1 U1729 ( .I(V84[16]), .ZN(n1629) );
  or2 U1730 ( .A1(n1744), .A2(n1629), .Z(n1526) );
  and2 U1731 ( .A1(n1527), .A2(n1526), .Z(n1531) );
  inv1 U1732 ( .I(V116[16]), .ZN(n1528) );
  or2 U1733 ( .A1(n1529), .A2(n1528), .Z(n1530) );
  and2 U1734 ( .A1(V84[5]), .A2(n876), .Z(n1535) );
  or2 U1735 ( .A1(n1753), .A2(n1607), .Z(n1532) );
  inv1 U1736 ( .I(n1532), .ZN(n1533) );
  or2 U1737 ( .A1(n1533), .A2(n883), .Z(n1534) );
  or2 U1738 ( .A1(n1534), .A2(n1535), .Z(n1536) );
  or2 U1739 ( .A1(n849), .A2(n1536), .Z(V197[16]) );
  or2 U1741 ( .A1(n1743), .A2(n1644), .Z(n1538) );
  inv1 U1743 ( .I(n1540), .ZN(n1543) );
  inv1 U1744 ( .I(n1541), .ZN(n1542) );
  or2 U1745 ( .A1(n1543), .A2(n1542), .Z(n1549) );
  and2 U1746 ( .A1(V84[6]), .A2(n875), .Z(n1547) );
  or2 U1747 ( .A1(n1750), .A2(n1621), .Z(n1544) );
  inv1 U1748 ( .I(n1544), .ZN(n1545) );
  or2 U1749 ( .A1(n1545), .A2(n881), .Z(n1546) );
  or2 U1750 ( .A1(n1546), .A2(n1547), .Z(n1548) );
  or2 U1751 ( .A1(n1549), .A2(n1548), .Z(V197[17]) );
  or2 U1753 ( .A1(n1744), .A2(n1659), .Z(n1551) );
  and2 U1754 ( .A1(n1552), .A2(n1551), .Z(n1553) );
  inv1 U1755 ( .I(n1553), .ZN(n1556) );
  inv1 U1756 ( .I(n1554), .ZN(n1555) );
  or2 U1757 ( .A1(n1556), .A2(n1555), .Z(n1561) );
  and2 U1758 ( .A1(V84[7]), .A2(n1741), .Z(n1559) );
  or2 U1759 ( .A1(n1753), .A2(n1636), .Z(n1557) );
  inv1 U1760 ( .I(n1557), .ZN(n1558) );
  or2 U1761 ( .A1(n1561), .A2(n1560), .Z(V197[18]) );
  or2 U1763 ( .A1(n1745), .A2(n1674), .Z(n1563) );
  inv1 U1765 ( .I(n1565), .ZN(n1568) );
  inv1 U1766 ( .I(n1566), .ZN(n1567) );
  or2 U1767 ( .A1(n1568), .A2(n1567), .Z(n1572) );
  and2 U1768 ( .A1(V84[8]), .A2(n876), .Z(n1570) );
  or2 U1769 ( .A1(n830), .A2(n881), .Z(n1569) );
  or2 U1770 ( .A1(n1569), .A2(n1570), .Z(n1571) );
  or2 U1771 ( .A1(n1572), .A2(n1571), .Z(V197[19]) );
  or2 U1773 ( .A1(n1743), .A2(n1689), .Z(n1574) );
  and2 U1774 ( .A1(n1575), .A2(n1574), .Z(n1576) );
  inv1 U1775 ( .I(n1576), .ZN(n1579) );
  inv1 U1776 ( .I(n1577), .ZN(n1578) );
  or2 U1777 ( .A1(n1579), .A2(n1578), .Z(n1585) );
  and2 U1778 ( .A1(V84[9]), .A2(n876), .Z(n1583) );
  or2 U1779 ( .A1(n1750), .A2(n1666), .Z(n1580) );
  inv1 U1780 ( .I(n1580), .ZN(n1581) );
  or2 U1781 ( .A1(n1581), .A2(n881), .Z(n1582) );
  or2 U1782 ( .A1(n1582), .A2(n1583), .Z(n1584) );
  or2 U1783 ( .A1(n1585), .A2(n1584), .Z(V197[20]) );
  or2 U1785 ( .A1(n1745), .A2(n1704), .Z(n1587) );
  inv1 U1787 ( .I(n1589), .ZN(n1592) );
  inv1 U1788 ( .I(n1590), .ZN(n1591) );
  or2 U1789 ( .A1(n1592), .A2(n1591), .Z(n1597) );
  or2 U1791 ( .A1(n1751), .A2(n1681), .Z(n1593) );
  inv1 U1792 ( .I(n1593), .ZN(n1594) );
  or2 U1793 ( .A1(n1597), .A2(n1596), .Z(V197[21]) );
  or2 U1795 ( .A1(n1745), .A2(n1719), .Z(n1599) );
  inv1 U1796 ( .I(n1601), .ZN(n1602) );
  or2 U1797 ( .A1(n823), .A2(n1602), .Z(n1606) );
  and2 U1798 ( .A1(V84[11]), .A2(n875), .Z(n1604) );
  or2 U1799 ( .A1(n809), .A2(n882), .Z(n1603) );
  or2 U1800 ( .A1(n1604), .A2(n1603), .Z(n1605) );
  or2 U1801 ( .A1(n1606), .A2(n1605), .Z(V197[22]) );
  or2 U1803 ( .A1(n1745), .A2(n1608), .Z(n1609) );
  inv1 U1805 ( .I(n1611), .ZN(n1614) );
  inv1 U1806 ( .I(n1612), .ZN(n1613) );
  or2 U1807 ( .A1(n1614), .A2(n1613), .Z(n1620) );
  and2 U1808 ( .A1(V84[12]), .A2(n876), .Z(n1618) );
  or2 U1809 ( .A1(n1750), .A2(n1711), .Z(n1615) );
  inv1 U1810 ( .I(n1615), .ZN(n1616) );
  or2 U1811 ( .A1(n1616), .A2(n883), .Z(n1617) );
  or2 U1812 ( .A1(n1617), .A2(n1618), .Z(n1619) );
  or2 U1813 ( .A1(n1620), .A2(n1619), .Z(V197[23]) );
  or2 U1814 ( .A1(n806), .A2(n1621), .Z(n1624) );
  or2 U1815 ( .A1(n1746), .A2(n1622), .Z(n1623) );
  and2 U1816 ( .A1(n1624), .A2(n1623), .Z(n1625) );
  inv1 U1818 ( .I(n1626), .ZN(n1627) );
  or2 U1819 ( .A1(n1628), .A2(n1627), .Z(n1635) );
  and2 U1820 ( .A1(V84[13]), .A2(n876), .Z(n1633) );
  or2 U1821 ( .A1(n1751), .A2(n1629), .Z(n1630) );
  inv1 U1822 ( .I(n1630), .ZN(n1631) );
  or2 U1823 ( .A1(n1631), .A2(n883), .Z(n1632) );
  or2 U1824 ( .A1(n1632), .A2(n1633), .Z(n1634) );
  or2 U1825 ( .A1(n1635), .A2(n1634), .Z(V197[24]) );
  or2 U1827 ( .A1(n1743), .A2(n1637), .Z(n1638) );
  inv1 U1830 ( .I(n1641), .ZN(n1642) );
  or2 U1831 ( .A1(n1643), .A2(n1642), .Z(n1650) );
  and2 U1832 ( .A1(V84[14]), .A2(n876), .Z(n1648) );
  or2 U1833 ( .A1(n1748), .A2(n1644), .Z(n1645) );
  inv1 U1834 ( .I(n1645), .ZN(n1646) );
  or2 U1835 ( .A1(n1646), .A2(n881), .Z(n1647) );
  or2 U1836 ( .A1(n1647), .A2(n1648), .Z(n1649) );
  or2 U1837 ( .A1(n1650), .A2(n1649), .Z(V197[25]) );
  or2 U1838 ( .A1(n803), .A2(n1651), .Z(n1654) );
  or2 U1839 ( .A1(n1746), .A2(n1652), .Z(n1653) );
  inv1 U1841 ( .I(n1655), .ZN(n1658) );
  inv1 U1842 ( .I(n1656), .ZN(n1657) );
  or2 U1843 ( .A1(n1658), .A2(n1657), .Z(n1665) );
  and2 U1844 ( .A1(V84[15]), .A2(n1740), .Z(n1663) );
  or2 U1845 ( .A1(n1750), .A2(n1659), .Z(n1660) );
  inv1 U1846 ( .I(n1660), .ZN(n1661) );
  or2 U1847 ( .A1(n1661), .A2(n882), .Z(n1662) );
  or2 U1848 ( .A1(n1662), .A2(n1663), .Z(n1664) );
  or2 U1849 ( .A1(n1665), .A2(n1664), .Z(V197[26]) );
  or2 U1850 ( .A1(n806), .A2(n1666), .Z(n1669) );
  or2 U1851 ( .A1(n1747), .A2(n1667), .Z(n1668) );
  and2 U1852 ( .A1(n1669), .A2(n1668), .Z(n1670) );
  inv1 U1854 ( .I(n1671), .ZN(n1672) );
  or2 U1855 ( .A1(n1673), .A2(n1672), .Z(n1680) );
  and2 U1856 ( .A1(V84[16]), .A2(n1740), .Z(n1678) );
  or2 U1857 ( .A1(n1752), .A2(n1674), .Z(n1675) );
  inv1 U1858 ( .I(n1675), .ZN(n1676) );
  or2 U1859 ( .A1(n1676), .A2(n883), .Z(n1677) );
  or2 U1860 ( .A1(n1677), .A2(n1678), .Z(n1679) );
  or2 U1861 ( .A1(n1680), .A2(n1679), .Z(V197[27]) );
  or2 U1862 ( .A1(n806), .A2(n1681), .Z(n1684) );
  or2 U1863 ( .A1(n1746), .A2(n1682), .Z(n1683) );
  and2 U1864 ( .A1(n1684), .A2(n1683), .Z(n1685) );
  inv1 U1866 ( .I(n1686), .ZN(n1687) );
  or2 U1867 ( .A1(n1688), .A2(n1687), .Z(n1695) );
  and2 U1868 ( .A1(V84[17]), .A2(n876), .Z(n1693) );
  or2 U1869 ( .A1(n1748), .A2(n1689), .Z(n1690) );
  inv1 U1870 ( .I(n1690), .ZN(n1691) );
  or2 U1871 ( .A1(n1691), .A2(n882), .Z(n1692) );
  or2 U1872 ( .A1(n1693), .A2(n1692), .Z(n1694) );
  or2 U1873 ( .A1(n1695), .A2(n1694), .Z(V197[28]) );
  or2 U1875 ( .A1(n1747), .A2(n1697), .Z(n1698) );
  and2 U1876 ( .A1(n1699), .A2(n1698), .Z(n1700) );
  inv1 U1877 ( .I(n1700), .ZN(n1703) );
  inv1 U1878 ( .I(n1701), .ZN(n1702) );
  or2 U1879 ( .A1(n1703), .A2(n1702), .Z(n1710) );
  and2 U1880 ( .A1(V84[18]), .A2(n876), .Z(n1708) );
  or2 U1881 ( .A1(n1748), .A2(n1704), .Z(n1705) );
  inv1 U1882 ( .I(n1705), .ZN(n1706) );
  or2 U1883 ( .A1(n1706), .A2(n881), .Z(n1707) );
  or2 U1884 ( .A1(n1707), .A2(n1708), .Z(n1709) );
  or2 U1885 ( .A1(n1710), .A2(n1709), .Z(V197[29]) );
  or2 U1886 ( .A1(n806), .A2(n1711), .Z(n1714) );
  or2 U1887 ( .A1(n1743), .A2(n1712), .Z(n1713) );
  and2 U1888 ( .A1(n1714), .A2(n1713), .Z(n1715) );
  inv1 U1890 ( .I(n1716), .ZN(n1717) );
  or2 U1891 ( .A1(n1718), .A2(n1717), .Z(n1725) );
  and2 U1892 ( .A1(V84[19]), .A2(n875), .Z(n1723) );
  or2 U1893 ( .A1(n1752), .A2(n1719), .Z(n1720) );
  inv1 U1894 ( .I(n1720), .ZN(n1721) );
  or2 U1895 ( .A1(n1721), .A2(n882), .Z(n1722) );
  or2 U1896 ( .A1(n1722), .A2(n1723), .Z(n1724) );
  or2 U1897 ( .A1(n1725), .A2(n1724), .Z(V197[30]) );
  and2 U1898 ( .A1(n874), .A2(V84[23]), .Z(n1728) );
  and2 U1899 ( .A1(V84[20]), .A2(n875), .Z(n1727) );
  or2 U1900 ( .A1(n1728), .A2(n1727), .Z(n1731) );
  and2 U1901 ( .A1(n800), .A2(V84[16]), .Z(n1730) );
  or2 U1902 ( .A1(n1731), .A2(n1730), .Z(n1737) );
  and2 U1903 ( .A1(n813), .A2(V84[31]), .Z(n1733) );
  or2 U1904 ( .A1(n1734), .A2(n1733), .Z(n1735) );
  or2 U1905 ( .A1(n881), .A2(n1735), .Z(n1736) );
  or2 U1906 ( .A1(n1737), .A2(n1736), .Z(V197[31]) );
  inv1 U856 ( .I(n1358), .ZN(n1740) );
  inv1 U857 ( .I(n1358), .ZN(n1741) );
  inv1f U859 ( .I(n868), .ZN(n871) );
  inv1 U861 ( .I(n1358), .ZN(n875) );
  or2 U862 ( .A1(n23), .A2(n1044), .Z(V143[0]) );
  or2 U863 ( .A1(n805), .A2(n1586), .Z(n1588) );
  and2f U870 ( .A1(n1588), .A2(n1587), .Z(n1589) );
  or2 U871 ( .A1(n802), .A2(n1537), .Z(n1539) );
  and2f U873 ( .A1(n1539), .A2(n1538), .Z(n1540) );
  and2f U878 ( .A1(n1639), .A2(n1638), .Z(n1640) );
  or2 U882 ( .A1(n801), .A2(n1636), .Z(n1639) );
  and2f U885 ( .A1(n1454), .A2(n1453), .Z(n1455) );
  or2 U887 ( .A1(n843), .A2(n1452), .Z(n1454) );
  and2f U888 ( .A1(n1045), .A2(V47[1]), .Z(n1035) );
  and2f U889 ( .A1(n1045), .A2(V47[8]), .Z(n1139) );
  or2 U890 ( .A1(n802), .A2(n1562), .Z(n1564) );
  and2f U891 ( .A1(n1564), .A2(n1563), .Z(n1565) );
  and2f U892 ( .A1(V84[5]), .A2(n1141), .Z(n1002) );
  and2f U893 ( .A1(V84[4]), .A2(n1141), .Z(n995) );
  and2f U900 ( .A1(V84[9]), .A2(n1141), .Z(n1036) );
  and2f U901 ( .A1(V47[5]), .A2(n1141), .Z(n1142) );
  and2f U902 ( .A1(n1063), .A2(n1032), .Z(n1033) );
  or2f U903 ( .A1(n1052), .A2(n1051), .Z(n1053) );
  or2f U904 ( .A1(n1061), .A2(n1060), .Z(n1062) );
  or2 U905 ( .A1(n835), .A2(V133[1]), .Z(n1088) );
  or2f U906 ( .A1(n1101), .A2(V133[6]), .Z(n835) );
  and2f U908 ( .A1(n1463), .A2(n1462), .Z(n1464) );
  inv1f U910 ( .I(n1726), .ZN(n837) );
  or2f U911 ( .A1(n1331), .A2(n1330), .Z(n1337) );
  inv1f U916 ( .I(n1092), .ZN(n865) );
  inv1 U917 ( .I(n386), .ZN(n1342) );
  or2 U918 ( .A1(n1140), .A2(n1055), .Z(n1057) );
  or2 U920 ( .A1(n1071), .A2(n1070), .Z(n1081) );
  or2 U922 ( .A1(n869), .A2(n1492), .Z(n1311) );
  inv1 U923 ( .I(V133[1]), .ZN(n778) );
  or2 U924 ( .A1(n949), .A2(n948), .Z(n1024) );
  and2 U925 ( .A1(n941), .A2(V133[1]), .Z(n807) );
  inv1 U926 ( .I(n780), .ZN(n946) );
  and2 U927 ( .A1(V15[1]), .A2(n1144), .Z(n974) );
  inv1 U928 ( .I(n868), .ZN(n870) );
  inv1 U929 ( .I(n800), .ZN(n802) );
  inv1 U930 ( .I(n813), .ZN(n1747) );
  inv1 U938 ( .I(V133[9]), .ZN(n1738) );
  or2 U939 ( .A1(n1140), .A2(n1025), .Z(n1027) );
  or2 U940 ( .A1(n1140), .A2(n1035), .Z(n1037) );
  or2 U941 ( .A1(n1140), .A2(n1046), .Z(n1048) );
  and2 U943 ( .A1(V47[3]), .A2(n866), .Z(n1108) );
  or2 U944 ( .A1(n869), .A2(n1226), .Z(n1119) );
  or2 U948 ( .A1(n869), .A2(n1352), .Z(n1154) );
  or2 U950 ( .A1(n869), .A2(n1390), .Z(n1187) );
  or2 U951 ( .A1(n869), .A2(n1452), .Z(n1258) );
  and2 U952 ( .A1(V47[16]), .A2(n867), .Z(n1330) );
  inv1 U953 ( .I(n1455), .ZN(n1456) );
  inv1 U954 ( .I(n1505), .ZN(n821) );
  and2 U955 ( .A1(V84[10]), .A2(n1740), .Z(n1595) );
  inv1 U957 ( .I(n1640), .ZN(n1643) );
  or2 U958 ( .A1(n1001), .A2(n1000), .Z(V142[1]) );
  and2 U960 ( .A1(n1063), .A2(n1021), .Z(n1023) );
  and2 U961 ( .A1(n1063), .A2(n1062), .Z(n1064) );
  and2 U962 ( .A1(n1081), .A2(n1080), .Z(n1087) );
  or2 U964 ( .A1(n1152), .A2(n1151), .Z(V150[0]) );
  inv1 U965 ( .I(n1314), .ZN(n1322) );
  inv1 U966 ( .I(n1444), .ZN(n1445) );
  and2f U967 ( .A1(n1423), .A2(n1422), .Z(n1424) );
  or2 U971 ( .A1(n843), .A2(n1421), .Z(n1423) );
  and2f U976 ( .A1(V47[4]), .A2(n855), .Z(n996) );
  inv1f U982 ( .I(n1625), .ZN(n1628) );
  inv1f U983 ( .I(n1670), .ZN(n1673) );
  inv1f U984 ( .I(n1685), .ZN(n1688) );
  inv1f U1042 ( .I(n1715), .ZN(n1718) );
  or2f U1061 ( .A1(n803), .A2(n1472), .Z(n1474) );
  inv1f U1062 ( .I(n1732), .ZN(n1742) );
  inv1f U1063 ( .I(n1742), .ZN(n1743) );
  inv1f U1064 ( .I(n1742), .ZN(n1744) );
  inv1f U1065 ( .I(n1742), .ZN(n1745) );
  inv1f U1066 ( .I(n813), .ZN(n1746) );
  inv1 U1069 ( .I(n1732), .ZN(n813) );
  inv1 U1071 ( .I(n874), .ZN(n1748) );
  inv1 U1072 ( .I(n874), .ZN(n1749) );
  inv1 U1073 ( .I(n874), .ZN(n1750) );
  inv1 U1074 ( .I(n837), .ZN(n1751) );
  inv1 U1077 ( .I(n837), .ZN(n1752) );
  inv1 U1078 ( .I(n837), .ZN(n1753) );
  inv1 U1079 ( .I(n861), .ZN(n863) );
  inv1 U1080 ( .I(n804), .ZN(n805) );
  inv1 U1087 ( .I(n861), .ZN(n864) );
  and2f U1088 ( .A1(n1610), .A2(n1609), .Z(n1611) );
  or2 U1102 ( .A1(n801), .A2(n1607), .Z(n1610) );
  inv1f U1105 ( .I(n842), .ZN(n843) );
  and2f U1114 ( .A1(n1654), .A2(n1653), .Z(n1655) );
  or2f U1122 ( .A1(n803), .A2(n1481), .Z(n1483) );
  or2f U1126 ( .A1(n803), .A2(n1573), .Z(n1575) );
  or2f U1127 ( .A1(n803), .A2(n1598), .Z(n1600) );
  or2f U1132 ( .A1(V133[2]), .A2(V133[6]), .Z(n938) );
  and2f U1134 ( .A1(n1063), .A2(n1013), .Z(n1015) );
  inv1f U1135 ( .I(n1393), .ZN(n1394) );
  or2f U1146 ( .A1(n844), .A2(n1352), .Z(n1354) );
  or2f U1153 ( .A1(n824), .A2(n853), .Z(n937) );
  or2f U1154 ( .A1(n942), .A2(V133[0]), .Z(n943) );
  and2f U1158 ( .A1(V47[2]), .A2(n855), .Z(n973) );
  or2f U1165 ( .A1(n1341), .A2(V133[2]), .Z(n1074) );
  and2f U1168 ( .A1(n1063), .A2(n992), .Z(n994) );
  inv1f U1169 ( .I(n785), .ZN(n834) );
  and2f U1170 ( .A1(n1344), .A2(n1343), .Z(n1345) );
  or2 U1177 ( .A1(n1098), .A2(n1357), .Z(n1092) );
  or2 U1178 ( .A1(n1098), .A2(n1351), .Z(n1097) );
  or2f U1180 ( .A1(n1098), .A2(n786), .Z(n1328) );
  inv1f U1186 ( .I(n880), .ZN(n879) );
  or2f U1190 ( .A1(n805), .A2(n1550), .Z(n1552) );
  or2f U1196 ( .A1(n805), .A2(n1696), .Z(n1699) );
  inv1f U1197 ( .I(n1332), .ZN(n861) );
  or2f U1206 ( .A1(n801), .A2(n1503), .Z(n1505) );
  or2f U1209 ( .A1(n1020), .A2(n1019), .Z(n1021) );
  inv1f U1211 ( .I(n781), .ZN(n1045) );
  or2f U1212 ( .A1(n782), .A2(n856), .Z(n781) );
  and2f U1216 ( .A1(n1348), .A2(n1347), .Z(n1349) );
  inv1f U1225 ( .I(n842), .ZN(n844) );
  and2f U1226 ( .A1(n1443), .A2(n1442), .Z(n1444) );
  or2f U1229 ( .A1(n843), .A2(n1379), .Z(n1381) );
  and2f U1231 ( .A1(n947), .A2(n786), .Z(n780) );
  or2f U1235 ( .A1(n843), .A2(n1410), .Z(n1412) );
  or2f U1237 ( .A1(n843), .A2(n1368), .Z(n1370) );
  or2f U1248 ( .A1(n843), .A2(n1401), .Z(n1403) );
  or2f U1258 ( .A1(n802), .A2(n1525), .Z(n1527) );
  or2f U1281 ( .A1(n802), .A2(n1492), .Z(n1494) );
  or2f U1283 ( .A1(n801), .A2(n1512), .Z(n1514) );
  or2f U1290 ( .A1(n1361), .A2(n832), .Z(n1362) );
  inv1f U1292 ( .I(n804), .ZN(n806) );
  inv1f U1337 ( .I(n832), .ZN(n1140) );
  or2f U1431 ( .A1(n946), .A2(n854), .Z(n832) );
  and2f U1499 ( .A1(n1340), .A2(n922), .Z(n786) );
  or2f U1506 ( .A1(n951), .A2(n950), .Z(n1357) );
  or2f U1524 ( .A1(n1341), .A2(n852), .Z(n1344) );
  or2f U1525 ( .A1(n1361), .A2(n786), .Z(n1732) );
  or2 U1532 ( .A1(n844), .A2(n1461), .Z(n1463) );
  inv1f U1533 ( .I(n880), .ZN(n878) );
  and2f U1535 ( .A1(n1360), .A2(n786), .Z(n857) );
  or2f U1536 ( .A1(n948), .A2(n834), .Z(n944) );
  inv1f U1539 ( .I(n1092), .ZN(n866) );
  and2f U1540 ( .A1(n824), .A2(n396), .Z(n77) );
  inv1f U1541 ( .I(n879), .ZN(n804) );
  inv1f U1542 ( .I(n879), .ZN(n842) );
  or2f U1543 ( .A1(n1078), .A2(n1077), .Z(n1090) );
  or2f U1549 ( .A1(n1076), .A2(n1075), .Z(n1077) );
  inv1f U1551 ( .I(n939), .ZN(n940) );
  or2f U1554 ( .A1(n938), .A2(V133[5]), .Z(n939) );
  inv1f U1558 ( .I(n1351), .ZN(n1144) );
  or2f U1570 ( .A1(n946), .A2(n945), .Z(n1351) );
  and2f U1586 ( .A1(n777), .A2(n778), .Z(n776) );
  and2f U1594 ( .A1(V133[5]), .A2(n776), .Z(n386) );
  and2f U1604 ( .A1(n1350), .A2(n1349), .Z(n775) );
  inv1f U1616 ( .I(n1726), .ZN(n874) );
  or2f U1619 ( .A1(n946), .A2(n854), .Z(n1360) );
  and2f U1641 ( .A1(V47[1]), .A2(n855), .Z(n960) );
  and2f U1642 ( .A1(V47[5]), .A2(n855), .Z(n1003) );
  or2f U1650 ( .A1(n781), .A2(n1098), .Z(n1332) );
  or2f U1653 ( .A1(V133[10]), .A2(n396), .Z(n1075) );
  and2f U1654 ( .A1(n1738), .A2(V133[7]), .Z(n396) );
  inv1f U1660 ( .I(V133[2]), .ZN(n853) );
  or2f U1663 ( .A1(n824), .A2(n853), .Z(n825) );
  or2f U1672 ( .A1(n937), .A2(n1072), .Z(n1340) );
  or2f U1682 ( .A1(n1024), .A2(n856), .Z(n950) );
  inv1f U1694 ( .I(n1357), .ZN(n1141) );
  inv1f U1706 ( .I(n1097), .ZN(n867) );
  and2f U1716 ( .A1(n941), .A2(V133[1]), .Z(n949) );
  or2f U1728 ( .A1(n940), .A2(V133[8]), .Z(n941) );
  or2f U1740 ( .A1(n775), .A2(n781), .Z(n1726) );
  or2f U1742 ( .A1(n775), .A2(n1357), .Z(n1358) );
  inv1f U1752 ( .I(n1729), .ZN(n880) );
  or2f U1762 ( .A1(n1361), .A2(n1351), .Z(n1729) );
  inv1f U1764 ( .I(V133[1]), .ZN(n824) );
  and2f U1772 ( .A1(n1350), .A2(n1349), .Z(n1361) );
  and2f U1784 ( .A1(n1345), .A2(n1346), .Z(n1350) );
  inv1f U1786 ( .I(n800), .ZN(n803) );
  inv1f U1790 ( .I(n878), .ZN(n800) );
  inv1f U1794 ( .I(n857), .ZN(n855) );
  or2f U1802 ( .A1(n945), .A2(n959), .Z(n854) );
  or2f U1804 ( .A1(n807), .A2(n944), .Z(n945) );
  or2f U1817 ( .A1(n1101), .A2(V133[6]), .Z(n1341) );
  or2f U1826 ( .A1(V133[9]), .A2(V133[4]), .Z(n1101) );
  inv1f U1828 ( .I(n1136), .ZN(n1098) );
  or2f U1829 ( .A1(n1090), .A2(n1089), .Z(n1136) );
  inv1f U1840 ( .I(n1328), .ZN(n868) );
endmodule

