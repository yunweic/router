
module k2 ( s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, 
        b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, 
        e, d, c, b, a, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, 
        x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, 
        f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0 );
  input s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0,
         a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e,
         d, c, b, a;
  output l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1,
         u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1,
         d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0;
  wire   n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n45, n50, n51, n52, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n68, n75, n76, n77, n78, n81, n85, n87, n91, n92, n93, n97, n98,
         n99, n100, n103, n105, n106, n108, n109, n112, n113, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n148, n149, n150, n151, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n171, n172, n174, n175, n176, n177, n178, n179, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n197, n198, n199, n200, n203, n204, n207, n208, n209,
         n210, n213, n214, n215, n216, n221, n223, n225, n226, n227, n228,
         n229, n230, n232, n233, n234, n237, n238, n239, n242, n243, n246,
         n247, n249, n250, n251, n252, n253, n254, n255, n256, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n276, n277, n278, n279, n281, n283, n284, n288, n289, n290,
         n294, n296, n297, n298, n299, n308, n309, n310, n311, n312, n313,
         n314, n317, n323, n325, n326, n327, n328, n329, n338, n343, n344,
         n346, n347, n348, n355, n356, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n375, n376, n382,
         n383, n384, n389, n390, n397, n398, n402, n404, n410, n419, n420,
         n421, n424, n425, n431, n451, n468, n473, n476, n483, n492, n493,
         n494, n495, n496, n497, n506, n507, n508, n509, n510, n511, n512,
         n516, n517, n518, n524, n525, n526, n527, n528, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n547, n548,
         n550, n551, n552, n553, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n570, n571, n572, n573, n575, n576, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n597, n602, n605, n606, n607, n608, n609, n610, n611, n616,
         n624, n625, n626, n630, n631, n632, n633, n634, n635, n636, n638,
         n640, n641, n642, n643, n644, n645, n646, n648, n649, n651, n652,
         n653, n656, n657, n664, n665, n669, n670, n671, n672, n674, n676,
         n686, n691, n692, n696, n697, n699, n700, n709, n714, n715, n716,
         n719, n722, n723, n725, n728, n732, n733, n734, n735, n736, n748,
         n749, n750, n751, n752, n753, n754, n755, n757, n768, n769, n770,
         n774, n777, n778, n781, n782, n784, n785, n786, n787, n788, n789,
         n790, n793, n796, n802, n803, n808, n809, n810, n832, n841, n842,
         n843, n844, n846, n847, n848, n849, n850, n851, n854, n861, n862,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1098, n1099, n1100,
         n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1162, n1163, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501;

  or2f U34 ( .A1(n97), .A2(n98), .Z(n75) );
  or2f U35 ( .A1(n99), .A2(n100), .Z(n98) );
  or2f U45 ( .A1(n117), .A2(n118), .Z(n116) );
  or2f U55 ( .A1(n134), .A2(n135), .Z(k1) );
  or2f U56 ( .A1(n136), .A2(n137), .Z(n135) );
  or2f U57 ( .A1(n138), .A2(n139), .Z(n137) );
  or2f U60 ( .A1(n143), .A2(n144), .Z(n120) );
  or2f U61 ( .A1(n145), .A2(n146), .Z(n144) );
  or2f U70 ( .A1(n161), .A2(n162), .Z(j1) );
  or2f U71 ( .A1(n163), .A2(n164), .Z(n162) );
  or2f U72 ( .A1(n165), .A2(n166), .Z(n164) );
  or2f U76 ( .A1(n1401), .A2(n1372), .Z(n169) );
  or2f U77 ( .A1(n171), .A2(n172), .Z(n1401) );
  or2f U84 ( .A1(n183), .A2(n184), .Z(i1) );
  or2f U92 ( .A1(n133), .A2(n68), .Z(n193) );
  or2f U97 ( .A1(n1353), .A2(n875), .Z(n199) );
  or2f U98 ( .A1(n203), .A2(n204), .Z(n197) );
  or2f U100 ( .A1(n207), .A2(n208), .Z(n183) );
  or2f U103 ( .A1(n1360), .A2(n213), .Z(n207) );
  or2f U104 ( .A1(n1395), .A2(n1366), .Z(n213) );
  or2f U112 ( .A1(n225), .A2(n226), .Z(n1395) );
  or2f U121 ( .A1(n237), .A2(n238), .Z(n78) );
  or2f U122 ( .A1(n191), .A2(n239), .Z(n238) );
  or2f U123 ( .A1(n1373), .A2(n1362), .Z(n239) );
  and2f U136 ( .A1(n256), .A2(n1431), .Z(n255) );
  or2f U137 ( .A1(n1380), .A2(n259), .Z(n256) );
  or2f U138 ( .A1(n260), .A2(n261), .Z(n259) );
  or2f U141 ( .A1(n265), .A2(n266), .Z(n264) );
  and2f U142 ( .A1(t), .A2(n267), .Z(n266) );
  or2f U143 ( .A1(n268), .A2(n269), .Z(n267) );
  and2f U144 ( .A1(u), .A2(n270), .Z(n269) );
  and2f U183 ( .A1(u), .A2(n326), .Z(n310) );
  or2f U184 ( .A1(n327), .A2(n328), .Z(n326) );
  and2f U185 ( .A1(v), .A2(n329), .Z(n328) );
  or2f U219 ( .A1(n363), .A2(n364), .Z(n139) );
  or2f U220 ( .A1(n365), .A2(n366), .Z(n364) );
  or2f U221 ( .A1(n234), .A2(n367), .Z(n366) );
  or2f U248 ( .A1(n1355), .A2(n402), .Z(n397) );
  and2f U251 ( .A1(a0), .A2(n404), .Z(n127) );
  and2f U271 ( .A1(n1386), .A2(n1384), .Z(n425) );
  or2f U360 ( .A1(n508), .A2(n509), .Z(n367) );
  or2f U361 ( .A1(n510), .A2(n511), .Z(n509) );
  or2f U362 ( .A1(n431), .A2(n512), .Z(n508) );
  or2f U363 ( .A1(n1359), .A2(n468), .Z(n512) );
  and2f U366 ( .A1(n517), .A2(n518), .Z(n516) );
  or2f U372 ( .A1(n527), .A2(n526), .Z(n99) );
  or2f U373 ( .A1(n528), .A2(n119), .Z(n527) );
  or2f U374 ( .A1(n187), .A2(n1435), .Z(n526) );
  or2f U380 ( .A1(n535), .A2(n536), .Z(n383) );
  or2f U381 ( .A1(n537), .A2(n538), .Z(n536) );
  and2f U388 ( .A1(n548), .A2(n1154), .Z(n547) );
  and2f U392 ( .A1(n551), .A2(n494), .Z(n537) );
  or2f U403 ( .A1(n559), .A2(n560), .Z(n535) );
  and2f U410 ( .A1(n565), .A2(n1357), .Z(n539) );
  or2f U430 ( .A1(n589), .A2(n588), .Z(n119) );
  or2f U431 ( .A1(n194), .A2(n590), .Z(n589) );
  and2f U454 ( .A1(x), .A2(n611), .Z(n106) );
  and2f U455 ( .A1(n611), .A2(w), .Z(n610) );
  and2f U456 ( .A1(b), .A2(n1361), .Z(n611) );
  or2f U472 ( .A1(n624), .A2(n625), .Z(n533) );
  or2f U481 ( .A1(n632), .A2(n633), .Z(n227) );
  or2f U482 ( .A1(n148), .A2(n573), .Z(n633) );
  or2f U484 ( .A1(n1403), .A2(n869), .Z(n634) );
  or2f U491 ( .A1(n640), .A2(n641), .Z(n590) );
  or2f U492 ( .A1(n642), .A2(n643), .Z(n641) );
  and2f U494 ( .A1(n390), .A2(n644), .Z(n642) );
  or2f U496 ( .A1(n646), .A2(n645), .Z(n640) );
  or2f U497 ( .A1(n648), .A2(n865), .Z(n646) );
  and2f U502 ( .A1(n635), .A2(n651), .Z(n645) );
  and2f U504 ( .A1(n1378), .A2(n1444), .Z(n635) );
  or2f U523 ( .A1(n669), .A2(n670), .Z(n572) );
  or2f U524 ( .A1(n671), .A2(n672), .Z(n670) );
  and2f U526 ( .A1(n674), .A2(n1376), .Z(n671) );
  or2f U546 ( .A1(n691), .A2(n692), .Z(n1402) );
  and2f U555 ( .A1(n1365), .A2(n700), .Z(n699) );
  or2f U580 ( .A1(n714), .A2(n715), .Z(n1409) );
  or2f U585 ( .A1(n1383), .A2(n1366), .Z(n714) );
  or2f U589 ( .A1(n561), .A2(n722), .Z(n203) );
  and2f U603 ( .A1(n733), .A2(n1386), .Z(n159) );
  or2f U604 ( .A1(n734), .A2(n735), .Z(n733) );
  and2f U605 ( .A1(d), .A2(n1384), .Z(n735) );
  and2f U606 ( .A1(w), .A2(n1382), .Z(n734) );
  or2f U619 ( .A1(n749), .A2(n750), .Z(n748) );
  or2f U620 ( .A1(n534), .A2(n585), .Z(n750) );
  or2f U621 ( .A1(n751), .A2(n752), .Z(n534) );
  or2f U622 ( .A1(n753), .A2(n754), .Z(n752) );
  or2f U623 ( .A1(n142), .A2(n510), .Z(n754) );
  or2f U624 ( .A1(n87), .A2(n755), .Z(n510) );
  and2f U627 ( .A1(n1468), .A2(n841), .Z(n757) );
  and2f U631 ( .A1(n518), .A2(n652), .Z(n87) );
  or2f U642 ( .A1(n768), .A2(n769), .Z(n751) );
  and2f U645 ( .A1(n278), .A2(n631), .Z(n770) );
  or2f U649 ( .A1(n1411), .A2(n58), .Z(n768) );
  or2f U656 ( .A1(n1372), .A2(n774), .Z(n585) );
  or2f U657 ( .A1(n242), .A2(n1373), .Z(n774) );
  and2f U660 ( .A1(n777), .A2(n778), .Z(n242) );
  or2f U667 ( .A1(n781), .A2(n782), .Z(n511) );
  or2f U668 ( .A1(n85), .A2(n81), .Z(n782) );
  and2f U669 ( .A1(w), .A2(n518), .Z(n81) );
  or2f U672 ( .A1(n221), .A2(n597), .Z(n781) );
  or2f U677 ( .A1(n784), .A2(n785), .Z(n194) );
  or2f U678 ( .A1(n786), .A2(n787), .Z(n785) );
  or2f U684 ( .A1(n676), .A2(n788), .Z(n784) );
  and2f U686 ( .A1(n1391), .A2(a0), .Z(n283) );
  and2f U688 ( .A1(r), .A2(n789), .Z(n676) );
  and2f U689 ( .A1(n1378), .A2(n1439), .Z(n789) );
  and2f U690 ( .A1(n1378), .A2(n790), .Z(n607) );
  and2f U785 ( .A1(a), .A2(n1384), .Z(n842) );
  and2f U789 ( .A1(n548), .A2(n525), .Z(n390) );
  and2f U802 ( .A1(n1476), .A2(n1425), .Z(n696) );
  and2f U817 ( .A1(n1390), .A2(u), .Z(n548) );
  and2f U822 ( .A1(n278), .A2(n421), .Z(n626) );
  and2f U838 ( .A1(n299), .A2(n525), .Z(n421) );
  and2f U839 ( .A1(t), .A2(d0), .Z(n525) );
  and2f U865 ( .A1(n1258), .A2(n1370), .Z(n861) );
  and2f U881 ( .A1(n876), .A2(d), .Z(n875) );
  buf0 U883 ( .I(n1412), .Z(u0) );
  buf0 U884 ( .I(n1411), .Z(w0) );
  buf0 U885 ( .I(n1410), .Z(x0) );
  buf0 U886 ( .I(n1409), .Z(y0) );
  buf0 U887 ( .I(n1408), .Z(b1) );
  buf0 U888 ( .I(n1407), .Z(c1) );
  buf0 U889 ( .I(n1406), .Z(h1) );
  buf0 U890 ( .I(n1405), .Z(n1) );
  buf0 U891 ( .I(n1404), .Z(o1) );
  buf0 U892 ( .I(n1403), .Z(q1) );
  buf0 U893 ( .I(n1350), .Z(r1) );
  buf0 U894 ( .I(n1402), .Z(t1) );
  buf0 U895 ( .I(n1401), .Z(u1) );
  buf0 U896 ( .I(n1400), .Z(v1) );
  buf0 U897 ( .I(n1399), .Z(x1) );
  buf0 U898 ( .I(n1398), .Z(y1) );
  buf0 U899 ( .I(n1397), .Z(z1) );
  buf0 U900 ( .I(n1396), .Z(c2) );
  buf0 U901 ( .I(n1395), .Z(g2) );
  buf0 U902 ( .I(n1394), .Z(i2) );
  buf0 U903 ( .I(n1393), .Z(k2) );
  buf0 U904 ( .I(n1350), .Z(l2) );
  or2 U905 ( .A1(n1280), .A2(n1478), .Z(n1173) );
  or2 U906 ( .A1(n1166), .A2(j), .Z(n938) );
  or2 U907 ( .A1(n1186), .A2(n1389), .Z(n1165) );
  inv1 U908 ( .I(n1166), .ZN(n1168) );
  and2f U909 ( .A1(e0), .A2(u), .Z(n899) );
  inv1f U910 ( .I(n899), .ZN(n1197) );
  or2 U911 ( .A1(n1489), .A2(n1441), .Z(n1085) );
  inv1 U912 ( .I(n1240), .ZN(n1241) );
  or2 U916 ( .A1(n1279), .A2(n1393), .Z(n1228) );
  and2 U917 ( .A1(n609), .A2(n1390), .Z(n664) );
  or2 U918 ( .A1(n1495), .A2(n1210), .Z(n1199) );
  or2 U919 ( .A1(n1495), .A2(f), .Z(n920) );
  or2 U920 ( .A1(n1390), .A2(n1431), .Z(n904) );
  inv1f U923 ( .I(e0), .ZN(n1390) );
  and2f U927 ( .A1(n1476), .A2(n1471), .Z(n851) );
  and2f U929 ( .A1(n626), .A2(n899), .Z(n901) );
  inv1f U936 ( .I(c0), .ZN(n1391) );
  inv1f U942 ( .I(n1204), .ZN(n1132) );
  or2f U943 ( .A1(n1132), .A2(n1391), .Z(n1033) );
  or2f U954 ( .A1(n1197), .A2(t), .Z(n1071) );
  inv1f U957 ( .I(n1133), .ZN(n1126) );
  or2f U963 ( .A1(n908), .A2(n907), .Z(n909) );
  and2f U964 ( .A1(n910), .A2(n909), .Z(n911) );
  or2f U965 ( .A1(n911), .A2(n579), .Z(n912) );
  or2f U966 ( .A1(n912), .A2(n582), .Z(n1255) );
  or2f U969 ( .A1(n1033), .A2(n913), .Z(n964) );
  or2f U970 ( .A1(n1491), .A2(n1431), .Z(n1240) );
  or2f U975 ( .A1(e0), .A2(u), .Z(n1008) );
  or2f U977 ( .A1(n1486), .A2(t), .Z(n1019) );
  or2f U978 ( .A1(n1019), .A2(n1008), .Z(n1042) );
  or2f U979 ( .A1(n1042), .A2(n1440), .Z(n1166) );
  or2f U983 ( .A1(n923), .A2(p0), .Z(n1005) );
  or2f U990 ( .A1(n1114), .A2(n1431), .Z(n921) );
  inv1f U991 ( .I(n921), .ZN(n45) );
  and2f U995 ( .A1(n1448), .A2(s), .Z(n925) );
  and2f U996 ( .A1(n925), .A2(n924), .Z(n1378) );
  or2f U1000 ( .A1(n1079), .A2(t), .Z(n1183) );
  or2f U1003 ( .A1(n980), .A2(n1068), .Z(n927) );
  or2f U1009 ( .A1(n1440), .A2(n936), .Z(n1049) );
  and2f U1016 ( .A1(n518), .A2(n1375), .Z(n597) );
  or2f U1018 ( .A1(n1198), .A2(c0), .Z(n1214) );
  and2f U1026 ( .A1(n934), .A2(n933), .Z(n1373) );
  or2f U1033 ( .A1(n941), .A2(n940), .Z(n942) );
  and2f U1045 ( .A1(n946), .A2(n1059), .Z(n247) );
  or2f U1053 ( .A1(n1183), .A2(d0), .Z(n1315) );
  or2f U1054 ( .A1(n953), .A2(n1315), .Z(n974) );
  or2f U1056 ( .A1(n974), .A2(n1190), .Z(n954) );
  and2f U1057 ( .A1(n955), .A2(n954), .Z(n956) );
  inv1f U1058 ( .I(n956), .ZN(n142) );
  or2f U1071 ( .A1(n748), .A2(n793), .Z(n969) );
  or2f U1077 ( .A1(n1467), .A2(n748), .Z(n1346) );
  inv1f U1078 ( .I(n1315), .ZN(n970) );
  and2f U1079 ( .A1(n970), .A2(n1148), .Z(n972) );
  or2f U1083 ( .A1(n973), .A2(n728), .Z(n1327) );
  or2f U1085 ( .A1(n974), .A2(f0), .Z(n975) );
  or2f U1086 ( .A1(n975), .A2(h0), .Z(n977) );
  and2f U1088 ( .A1(n977), .A2(n976), .Z(n978) );
  or2f U1090 ( .A1(n978), .A2(n1004), .Z(n979) );
  or2f U1101 ( .A1(n987), .A2(n1214), .Z(n988) );
  inv1f U1109 ( .I(n1074), .ZN(n1365) );
  or2f U1111 ( .A1(n991), .A2(n179), .Z(n691) );
  inv1f U1113 ( .I(n992), .ZN(n994) );
  or2f U1131 ( .A1(n1445), .A2(n1374), .Z(n644) );
  inv1f U1133 ( .I(n1214), .ZN(n1047) );
  and2f U1134 ( .A1(n1001), .A2(n1047), .Z(n643) );
  or2f U1136 ( .A1(n1002), .A2(n1441), .Z(n1003) );
  inv1f U1137 ( .I(n1003), .ZN(n156) );
  or2f U1138 ( .A1(n156), .A2(n636), .Z(n1403) );
  and2f U1142 ( .A1(n1204), .A2(n525), .Z(n1007) );
  and2f U1143 ( .A1(n1007), .A2(n1059), .Z(n1361) );
  or2f U1146 ( .A1(n1141), .A2(n591), .Z(n588) );
  or2f U1152 ( .A1(n602), .A2(n1405), .Z(n1016) );
  or2f U1156 ( .A1(n1404), .A2(n1014), .Z(n1015) );
  or2f U1157 ( .A1(n1016), .A2(n1015), .Z(n371) );
  or2f U1158 ( .A1(n121), .A2(n371), .Z(n228) );
  or2f U1169 ( .A1(n1385), .A2(n228), .Z(n1027) );
  or2f U1172 ( .A1(n1029), .A2(n1138), .Z(n1030) );
  or2f U1173 ( .A1(n1031), .A2(n1030), .Z(n1266) );
  or2f U1175 ( .A1(n1034), .A2(n1033), .Z(n1035) );
  or2f U1177 ( .A1(n1266), .A2(n1359), .Z(n1038) );
  or2f U1179 ( .A1(n1038), .A2(n1037), .Z(n583) );
  or2f U1185 ( .A1(n1077), .A2(f), .Z(n1044) );
  or2f U1187 ( .A1(c0), .A2(b0), .Z(n1045) );
  or2f U1188 ( .A1(n1045), .A2(d0), .Z(n1046) );
  or2f U1203 ( .A1(n1056), .A2(n1055), .Z(n1057) );
  and2f U1204 ( .A1(n1210), .A2(n1057), .Z(n1058) );
  and2f U1209 ( .A1(n1063), .A2(n1062), .Z(n1065) );
  or2f U1210 ( .A1(n1065), .A2(n1064), .Z(n1066) );
  or2f U1211 ( .A1(n1066), .A2(n516), .Z(n468) );
  or2f U1225 ( .A1(n1077), .A2(n1142), .Z(n1076) );
  and2f U1245 ( .A1(n1210), .A2(n1089), .Z(n1091) );
  and2f U1251 ( .A1(n1210), .A2(n1095), .Z(n327) );
  and2f U1266 ( .A1(n1117), .A2(n1107), .Z(n268) );
  or2f U1279 ( .A1(n1120), .A2(n308), .Z(n1121) );
  and2f U1282 ( .A1(n1458), .A2(n1123), .Z(n1124) );
  and2f U1289 ( .A1(n1129), .A2(n686), .Z(n1130) );
  and2f U1290 ( .A1(n1131), .A2(n1130), .Z(n182) );
  or2f U1294 ( .A1(n1402), .A2(n1475), .Z(n1135) );
  or2f U1295 ( .A1(n182), .A2(n1135), .Z(n62) );
  or2f U1300 ( .A1(n1138), .A2(n1268), .Z(n1139) );
  or2f U1301 ( .A1(n1140), .A2(n1139), .Z(n166) );
  or2f U1303 ( .A1(n1143), .A2(n1214), .Z(n1144) );
  inv1f U1304 ( .I(n1144), .ZN(n1211) );
  or2f U1308 ( .A1(n1232), .A2(n1387), .Z(n204) );
  and2f U1309 ( .A1(d), .A2(n1148), .Z(n1149) );
  or2f U1310 ( .A1(n1149), .A2(n1382), .Z(n1318) );
  and2f U1312 ( .A1(n1318), .A2(n1150), .Z(n200) );
  or2f U1321 ( .A1(n1166), .A2(n1154), .Z(n1155) );
  or2f U1334 ( .A1(n157), .A2(n1496), .Z(n1194) );
  or2f U1335 ( .A1(n151), .A2(n1194), .Z(n1172) );
  or2f U1340 ( .A1(n1172), .A2(n1171), .Z(n1280) );
  or2f U1347 ( .A1(n1301), .A2(n1178), .Z(n1179) );
  or2f U1360 ( .A1(n106), .A2(n75), .Z(n1196) );
  or2f U1362 ( .A1(n1196), .A2(n1195), .Z(n93) );
  or2f U1374 ( .A1(n1212), .A2(n1211), .Z(n1213) );
  or2f U1375 ( .A1(n1213), .A2(n1371), .Z(n1223) );
  or2f U1377 ( .A1(n1215), .A2(n1214), .Z(n1216) );
  or2f U1380 ( .A1(n1230), .A2(n1218), .Z(n1221) );
  or2f U1383 ( .A1(n1223), .A2(n1222), .Z(n1224) );
  and2f U1384 ( .A1(z), .A2(n1224), .Z(n1225) );
  and2f U1385 ( .A1(n1226), .A2(n1225), .Z(n1227) );
  and2f U1390 ( .A1(n1392), .A2(n861), .Z(n1234) );
  or2f U1391 ( .A1(n873), .A2(n1232), .Z(n1233) );
  or2f U1392 ( .A1(n1234), .A2(n1233), .Z(n1253) );
  and2f U1394 ( .A1(n1258), .A2(n1375), .Z(n1236) );
  or2f U1395 ( .A1(n1237), .A2(n1236), .Z(n1251) );
  and2f U1397 ( .A1(n1241), .A2(n1374), .Z(n1242) );
  and2f U1398 ( .A1(n1243), .A2(n1242), .Z(n1249) );
  or2f U1402 ( .A1(n1249), .A2(n1394), .Z(n1250) );
  or2f U1403 ( .A1(n1251), .A2(n1250), .Z(n1252) );
  or2f U1404 ( .A1(n1253), .A2(n1252), .Z(n1310) );
  or2f U1405 ( .A1(n1254), .A2(n1310), .Z(n1257) );
  or2f U1407 ( .A1(n1257), .A2(n1256), .Z(n1408) );
  or2f U1408 ( .A1(n1408), .A2(n578), .Z(n1264) );
  or2f U1411 ( .A1(n1260), .A2(n572), .Z(n1311) );
  or2f U1412 ( .A1(n1311), .A2(n1358), .Z(n1262) );
  or2f U1413 ( .A1(n1262), .A2(n1261), .Z(n1263) );
  or2f U1414 ( .A1(n1264), .A2(n1263), .Z(n1333) );
  or2f U1419 ( .A1(n1267), .A2(n1266), .Z(n1271) );
  or2f U1422 ( .A1(n1271), .A2(n1270), .Z(n1406) );
  or2f U1423 ( .A1(n75), .A2(n76), .Z(n1274) );
  or2f U1426 ( .A1(n1274), .A2(n1273), .Z(n1299) );
  or2f U1430 ( .A1(n1227), .A2(n1488), .Z(n1283) );
  or2f U1431 ( .A1(n468), .A2(n149), .Z(n1281) );
  or2f U1432 ( .A1(n1281), .A2(n1280), .Z(n1282) );
  or2f U1433 ( .A1(n1283), .A2(n1282), .Z(n1294) );
  or2f U1441 ( .A1(n1294), .A2(n1293), .Z(n1305) );
  or2f U1444 ( .A1(n1305), .A2(n1450), .Z(n1298) );
  or2f U1445 ( .A1(n1299), .A2(n1298), .Z(n1300) );
  or2f U1446 ( .A1(n1300), .A2(n1406), .Z(p1) );
  or2f U1453 ( .A1(n1305), .A2(n1462), .Z(n1308) );
  or2f U1454 ( .A1(n1309), .A2(n1308), .Z(n1400) );
  or2f U1458 ( .A1(n633), .A2(n1477), .Z(n1314) );
  or2f U1459 ( .A1(n1314), .A2(n533), .Z(n1324) );
  or2f U1465 ( .A1(n1324), .A2(n1323), .Z(n1332) );
  or2f U1471 ( .A1(n1332), .A2(n1331), .Z(n1334) );
  or2f U1472 ( .A1(n1333), .A2(n1334), .Z(n1396) );
  or2f U1483 ( .A1(n1345), .A2(n1344), .Z(n1347) );
  or2f U1484 ( .A1(n1346), .A2(n1347), .Z(n1348) );
  or2f U1485 ( .A1(n1348), .A2(n1396), .Z(n1349) );
  or2f U1486 ( .A1(n1349), .A2(n1400), .Z(e2) );
  inv1 U856 ( .I(1'b1), .ZN(v0) );
  inv1 U858 ( .I(1'b1), .ZN(j2) );
  or2f U860 ( .A1(n872), .A2(n868), .Z(n431) );
  or2f U861 ( .A1(n1098), .A2(n1434), .Z(n314) );
  inv1f U862 ( .I(n899), .ZN(n1495) );
  inv1f U863 ( .I(f), .ZN(n1142) );
  or2f U864 ( .A1(n1094), .A2(n1093), .Z(n329) );
  and2f U866 ( .A1(n1238), .A2(n1092), .Z(n1093) );
  inv1f U867 ( .I(n1023), .ZN(n1384) );
  or2f U868 ( .A1(n1033), .A2(n1201), .Z(n1023) );
  and2 U869 ( .A1(w), .A2(n1108), .Z(n1105) );
  or2 U870 ( .A1(n283), .A2(n284), .Z(n281) );
  or2 U871 ( .A1(n1091), .A2(n1090), .Z(n1092) );
  and2 U872 ( .A1(n949), .A2(n948), .Z(n246) );
  and2 U873 ( .A1(t), .A2(n314), .Z(n313) );
  inv1 U874 ( .I(n942), .ZN(n1371) );
  or2 U875 ( .A1(n1170), .A2(n1169), .Z(n1171) );
  or2 U876 ( .A1(n149), .A2(n150), .Z(n143) );
  and2 U877 ( .A1(n1126), .A2(n1125), .Z(n1127) );
  inv1 U878 ( .I(n985), .ZN(n1367) );
  and2 U879 ( .A1(n874), .A2(n1043), .Z(n873) );
  inv1 U880 ( .I(n1077), .ZN(n876) );
  or2 U882 ( .A1(n581), .A2(n1255), .Z(n1256) );
  and2 U913 ( .A1(n696), .A2(n697), .Z(n179) );
  or2 U914 ( .A1(n397), .A2(n398), .Z(n65) );
  or2 U915 ( .A1(n1354), .A2(n91), .Z(n398) );
  and2 U921 ( .A1(n1122), .A2(n1121), .Z(n254) );
  or2 U922 ( .A1(v), .A2(c0), .Z(n1423) );
  or2 U924 ( .A1(v), .A2(s), .Z(n1424) );
  inv1f U925 ( .I(n1424), .ZN(n1204) );
  inv1 U926 ( .I(s), .ZN(n1108) );
  or2 U928 ( .A1(n1068), .A2(n1446), .Z(n1077) );
  or2 U930 ( .A1(n1068), .A2(n1154), .Z(n985) );
  or2 U931 ( .A1(n1423), .A2(s), .Z(n1068) );
  inv1f U932 ( .I(n1434), .ZN(n1096) );
  and2 U933 ( .A1(n547), .A2(n1204), .Z(n1056) );
  and2 U934 ( .A1(n757), .A2(n548), .Z(n949) );
  and2f U935 ( .A1(n539), .A2(n540), .Z(n538) );
  or2f U937 ( .A1(n528), .A2(n1363), .Z(n148) );
  or2f U938 ( .A1(n246), .A2(n247), .Z(n755) );
  and2f U939 ( .A1(n262), .A2(n263), .Z(n261) );
  or2f U940 ( .A1(n1155), .A2(f0), .Z(n1191) );
  and2f U941 ( .A1(n631), .A2(a), .Z(n850) );
  inv1f U944 ( .I(d0), .ZN(n1486) );
  and2f U945 ( .A1(s), .A2(n1391), .Z(n1089) );
  and2f U946 ( .A1(n309), .A2(n1431), .Z(n308) );
  or2f U947 ( .A1(n1441), .A2(n960), .Z(n941) );
  inv1f U948 ( .I(n1471), .ZN(n960) );
  or2f U949 ( .A1(n1133), .A2(n1182), .Z(n1074) );
  and2f U950 ( .A1(a0), .A2(n841), .Z(n317) );
  and2f U951 ( .A1(n299), .A2(c0), .Z(n841) );
  and2 U952 ( .A1(n317), .A2(n1471), .Z(n946) );
  and2 U953 ( .A1(n1108), .A2(n1442), .Z(n1090) );
  or2 U955 ( .A1(w), .A2(z), .Z(n284) );
  inv1 U956 ( .I(n1484), .ZN(n1483) );
  inv1 U958 ( .I(f0), .ZN(n1485) );
  and2 U959 ( .A1(n1458), .A2(g), .Z(n1150) );
  and2 U960 ( .A1(c0), .A2(n770), .Z(n209) );
  inv1 U961 ( .I(n1036), .ZN(n1362) );
  and2 U962 ( .A1(n1479), .A2(n1012), .Z(n1014) );
  inv1 U967 ( .I(n1046), .ZN(n1357) );
  and2 U968 ( .A1(n1210), .A2(n1209), .Z(n1212) );
  inv1 U971 ( .I(n1217), .ZN(n1218) );
  inv1 U972 ( .I(n1219), .ZN(n1220) );
  or2 U973 ( .A1(n1370), .A2(w), .Z(n700) );
  and2 U974 ( .A1(n686), .A2(n609), .Z(n1123) );
  inv1 U976 ( .I(c0), .ZN(n1443) );
  inv1 U980 ( .I(n1033), .ZN(n1148) );
  or2 U981 ( .A1(n1111), .A2(n288), .Z(n1112) );
  and2 U982 ( .A1(u), .A2(n289), .Z(n288) );
  and2 U984 ( .A1(b), .A2(n657), .Z(n528) );
  or2 U985 ( .A1(n1183), .A2(n1182), .Z(n1219) );
  inv1 U986 ( .I(n1492), .ZN(n1494) );
  and2 U987 ( .A1(n1287), .A2(n1286), .Z(n1291) );
  or2 U988 ( .A1(l), .A2(n1081), .Z(n929) );
  and2 U989 ( .A1(n1204), .A2(n1442), .Z(n1376) );
  and2 U992 ( .A1(n1316), .A2(n1367), .Z(n991) );
  inv1 U993 ( .I(n1035), .ZN(n1359) );
  inv1 U994 ( .I(n1231), .ZN(n1370) );
  inv1 U997 ( .I(a), .ZN(n1431) );
  inv1 U998 ( .I(n932), .ZN(n778) );
  or2 U999 ( .A1(n372), .A2(n373), .Z(n363) );
  or2 U1001 ( .A1(n106), .A2(n610), .Z(n121) );
  or2 U1002 ( .A1(n78), .A2(n249), .Z(n1140) );
  or2 U1004 ( .A1(n197), .A2(n198), .Z(n174) );
  or2 U1005 ( .A1(n1369), .A2(n209), .Z(n769) );
  or2 U1006 ( .A1(n1362), .A2(n141), .Z(n625) );
  or2 U1007 ( .A1(n271), .A2(n272), .Z(n270) );
  and2 U1008 ( .A1(n518), .A2(n616), .Z(n868) );
  inv1 U1010 ( .I(n1165), .ZN(n1170) );
  and2 U1011 ( .A1(n1157), .A2(n1302), .Z(n151) );
  or2 U1012 ( .A1(n1191), .A2(n1162), .Z(n1163) );
  inv1 U1013 ( .I(n864), .ZN(n149) );
  and2 U1014 ( .A1(n1179), .A2(n1181), .Z(n864) );
  and2 U1015 ( .A1(n1476), .A2(n283), .Z(n686) );
  and2 U1017 ( .A1(n283), .A2(n1364), .Z(n672) );
  inv1 U1019 ( .I(n964), .ZN(n1382) );
  inv1 U1020 ( .I(n1301), .ZN(n1302) );
  and2 U1021 ( .A1(n605), .A2(n606), .Z(n602) );
  and2 U1022 ( .A1(a0), .A2(n1371), .Z(n59) );
  and2 U1023 ( .A1(n1083), .A2(n1376), .Z(n787) );
  inv1 U1024 ( .I(n927), .ZN(n786) );
  and2 U1025 ( .A1(n1479), .A2(n926), .Z(n788) );
  and2 U1027 ( .A1(n635), .A2(n517), .Z(n869) );
  or2 U1028 ( .A1(n371), .A2(n119), .Z(n365) );
  or2 U1029 ( .A1(n375), .A2(n1360), .Z(n372) );
  inv1 U1030 ( .I(x), .ZN(n1154) );
  inv1 U1031 ( .I(n1159), .ZN(n157) );
  or2 U1032 ( .A1(n1158), .A2(n1183), .Z(n1159) );
  or2 U1034 ( .A1(n242), .A2(n243), .Z(n237) );
  or2 U1035 ( .A1(n1221), .A2(n1220), .Z(n1222) );
  or2 U1036 ( .A1(n1124), .A2(n699), .Z(n1454) );
  and2 U1037 ( .A1(n548), .A2(n851), .Z(n631) );
  and2 U1038 ( .A1(n972), .A2(n971), .Z(n722) );
  inv1 U1039 ( .I(n914), .ZN(n1232) );
  and2 U1040 ( .A1(n1434), .A2(n810), .Z(n865) );
  inv1 U1041 ( .I(n979), .ZN(n983) );
  inv1 U1042 ( .I(d0), .ZN(n1472) );
  or2 U1043 ( .A1(n310), .A2(n311), .Z(n309) );
  and2 U1044 ( .A1(d0), .A2(n264), .Z(n262) );
  inv1 U1046 ( .I(n1076), .ZN(n1353) );
  and2 U1047 ( .A1(n1370), .A2(n1371), .Z(n55) );
  or2 U1048 ( .A1(n59), .A2(n55), .Z(n1411) );
  inv1 U1049 ( .I(n1041), .ZN(n1358) );
  or2 U1050 ( .A1(n141), .A2(n169), .Z(n77) );
  or2 U1051 ( .A1(n120), .A2(n140), .Z(n136) );
  inv1 U1052 ( .I(n1292), .ZN(n1293) );
  and2 U1055 ( .A1(n1291), .A2(n1290), .Z(n1292) );
  and2 U1059 ( .A1(n635), .A2(n638), .Z(n636) );
  or2 U1060 ( .A1(n994), .A2(n993), .Z(n692) );
  or2 U1061 ( .A1(n1259), .A2(n861), .Z(n1260) );
  or2 U1062 ( .A1(n990), .A2(n716), .Z(n715) );
  and2 U1063 ( .A1(b0), .A2(n696), .Z(n591) );
  or2 U1064 ( .A1(n918), .A2(n1391), .Z(n902) );
  and2 U1065 ( .A1(n850), .A2(n296), .Z(n561) );
  or2 U1066 ( .A1(n214), .A2(n383), .Z(n382) );
  or2 U1067 ( .A1(n968), .A2(n793), .Z(n1467) );
  and2 U1068 ( .A1(n901), .A2(n900), .Z(n1387) );
  or2 U1069 ( .A1(n1247), .A2(n1246), .Z(n1248) );
  or2 U1070 ( .A1(n1265), .A2(n1407), .Z(z0) );
  or2 U1072 ( .A1(n583), .A2(n584), .Z(d1) );
  or2 U1073 ( .A1(n361), .A2(n362), .Z(f1) );
  or2 U1074 ( .A1(n139), .A2(n165), .Z(n362) );
  or2 U1075 ( .A1(n232), .A2(n233), .Z(g1) );
  or2 U1076 ( .A1(n234), .A2(n166), .Z(n233) );
  or2 U1080 ( .A1(n185), .A2(n186), .Z(n184) );
  or2 U1081 ( .A1(n92), .A2(n93), .Z(m1) );
  or2 U1082 ( .A1(n60), .A2(n61), .Z(s1) );
  or2 U1084 ( .A1(n1229), .A2(n1228), .Z(n60) );
  or2 U1087 ( .A1(n530), .A2(n531), .Z(d2) );
  or2 U1089 ( .A1(n254), .A2(n255), .Z(n253) );
  inv1 U1091 ( .I(n1048), .ZN(n1425) );
  or2 U1092 ( .A1(n1402), .A2(n1475), .Z(n1426) );
  or2 U1093 ( .A1(n1426), .A2(n1427), .Z(n100) );
  or2 U1094 ( .A1(n1351), .A2(n182), .Z(n1427) );
  inv1 U1095 ( .I(n1048), .ZN(n1386) );
  and2 U1096 ( .A1(n1386), .A2(n1376), .Z(n993) );
  and2 U1097 ( .A1(n1377), .A2(n1386), .Z(n404) );
  and2 U1098 ( .A1(n649), .A2(n1432), .Z(n1469) );
  or2 U1099 ( .A1(n1061), .A2(n1445), .Z(n1062) );
  inv1f U1100 ( .I(n1049), .ZN(n1445) );
  or2f U1102 ( .A1(n1441), .A2(n1431), .Z(n1470) );
  inv1 U1103 ( .I(n1481), .ZN(n299) );
  inv1 U1104 ( .I(a), .ZN(n1244) );
  or2 U1105 ( .A1(n1245), .A2(n1244), .Z(n1490) );
  or2f U1106 ( .A1(f), .A2(p), .Z(n1245) );
  and2 U1107 ( .A1(s), .A2(v), .Z(n1428) );
  inv1f U1108 ( .I(n1428), .ZN(n1198) );
  inv1 U1110 ( .I(v), .ZN(n550) );
  or2 U1112 ( .A1(n1180), .A2(n1198), .Z(n1181) );
  or2 U1114 ( .A1(n969), .A2(n1498), .Z(n1429) );
  or2 U1115 ( .A1(n1429), .A2(n1430), .Z(b2) );
  or2 U1116 ( .A1(n725), .A2(n1026), .Z(n1430) );
  and2 U1117 ( .A1(n1316), .A2(n1047), .Z(n1050) );
  inv1 U1118 ( .I(n1198), .ZN(n1374) );
  or2 U1119 ( .A1(n1080), .A2(n1198), .Z(n1217) );
  or2 U1120 ( .A1(n1215), .A2(n1214), .Z(n1459) );
  inv1 U1121 ( .I(n1019), .ZN(n924) );
  and2f U1122 ( .A1(e0), .A2(n653), .Z(n518) );
  and2 U1123 ( .A1(v), .A2(n1378), .Z(n653) );
  inv1 U1124 ( .I(n1040), .ZN(n1364) );
  or2 U1125 ( .A1(n1040), .A2(n1231), .Z(n1041) );
  or2f U1126 ( .A1(n1008), .A2(n996), .Z(n1040) );
  and2f U1127 ( .A1(n1433), .A2(v), .Z(n1432) );
  inv1f U1128 ( .I(s), .ZN(n1433) );
  and2 U1129 ( .A1(n421), .A2(c0), .Z(n606) );
  and2f U1130 ( .A1(n283), .A2(n421), .Z(n926) );
  inv1 U1132 ( .I(n1481), .ZN(n1476) );
  or2f U1135 ( .A1(n227), .A2(n228), .Z(n226) );
  or2f U1139 ( .A1(n1315), .A2(n1068), .Z(n992) );
  or2f U1140 ( .A1(n1315), .A2(n1431), .Z(n987) );
  and2f U1141 ( .A1(n1432), .A2(c0), .Z(n1434) );
  or2 U1144 ( .A1(n1096), .A2(n1201), .Z(n1158) );
  or2 U1145 ( .A1(n1403), .A2(n209), .Z(n1435) );
  inv1 U1147 ( .I(n1436), .ZN(n187) );
  or2 U1148 ( .A1(n1078), .A2(n476), .Z(n1436) );
  and2 U1149 ( .A1(n317), .A2(n1117), .Z(n1098) );
  or2 U1150 ( .A1(n1214), .A2(n980), .Z(n930) );
  or2f U1151 ( .A1(n1183), .A2(n1472), .Z(n980) );
  or2f U1153 ( .A1(n1343), .A2(n382), .Z(n1345) );
  or2f U1154 ( .A1(n916), .A2(n915), .Z(n923) );
  or2 U1155 ( .A1(n383), .A2(n532), .Z(n531) );
  and2f U1159 ( .A1(n924), .A2(n548), .Z(n1437) );
  inv1f U1160 ( .I(n1437), .ZN(n1032) );
  inv1 U1161 ( .I(n548), .ZN(n986) );
  and2 U1162 ( .A1(r), .A2(n789), .Z(n1438) );
  and2 U1163 ( .A1(n1390), .A2(n790), .Z(n1439) );
  and2 U1164 ( .A1(n1438), .A2(a), .Z(n669) );
  and2 U1165 ( .A1(n607), .A2(n608), .Z(n1405) );
  inv1 U1166 ( .I(n1432), .ZN(n1441) );
  inv1f U1167 ( .I(n1432), .ZN(n1440) );
  and2f U1168 ( .A1(n1443), .A2(w), .Z(n1442) );
  inv1f U1170 ( .I(n1442), .ZN(n936) );
  inv1 U1171 ( .I(w), .ZN(n1201) );
  or2 U1174 ( .A1(n936), .A2(j), .Z(n915) );
  or2 U1176 ( .A1(n1197), .A2(t), .Z(n1456) );
  or2 U1178 ( .A1(n1049), .A2(n1048), .Z(n1246) );
  and2 U1180 ( .A1(u), .A2(n1432), .Z(n1209) );
  and2 U1181 ( .A1(n656), .A2(n1432), .Z(n1061) );
  and2 U1182 ( .A1(v), .A2(n1390), .Z(n1444) );
  or2 U1183 ( .A1(n1019), .A2(n1008), .Z(n1446) );
  or2 U1184 ( .A1(n923), .A2(n1447), .Z(n955) );
  or2 U1186 ( .A1(n1500), .A2(n950), .Z(n1447) );
  or2f U1189 ( .A1(n1071), .A2(d0), .Z(n1489) );
  and2f U1190 ( .A1(n1449), .A2(u), .Z(n1448) );
  inv1f U1191 ( .I(c0), .ZN(n1449) );
  or2 U1192 ( .A1(n1491), .A2(n1142), .Z(n1143) );
  or2f U1193 ( .A1(n590), .A2(n634), .Z(n573) );
  or2 U1194 ( .A1(n1297), .A2(n1501), .Z(n1450) );
  and2 U1195 ( .A1(n1226), .A2(n1225), .Z(n1451) );
  inv1 U1196 ( .I(n1453), .ZN(n1452) );
  inv1 U1197 ( .I(n1445), .ZN(n1453) );
  or2f U1198 ( .A1(n1454), .A2(n1455), .Z(n1475) );
  or2 U1199 ( .A1(n192), .A2(n1127), .Z(n1455) );
  or2f U1200 ( .A1(n1456), .A2(n1457), .Z(n1215) );
  or2f U1201 ( .A1(n1490), .A2(d0), .Z(n1457) );
  inv1f U1202 ( .I(n1489), .ZN(n1458) );
  or2 U1205 ( .A1(n1127), .A2(n168), .Z(n1128) );
  or2 U1206 ( .A1(n1124), .A2(n699), .Z(n168) );
  inv1f U1207 ( .I(n1489), .ZN(n1316) );
  or2 U1208 ( .A1(n1458), .A2(n1126), .Z(n1129) );
  and2 U1212 ( .A1(l), .A2(n1316), .Z(n908) );
  or2 U1213 ( .A1(n1128), .A2(n1402), .Z(n124) );
  or2 U1214 ( .A1(n1049), .A2(n952), .Z(n953) );
  or2f U1215 ( .A1(n983), .A2(n982), .Z(n1460) );
  or2f U1216 ( .A1(n1460), .A2(n1461), .Z(n1138) );
  or2f U1217 ( .A1(n1028), .A2(n1027), .Z(n1461) );
  or2 U1218 ( .A1(n1027), .A2(n1026), .Z(n1344) );
  or2 U1219 ( .A1(n983), .A2(n982), .Z(n1026) );
  or2f U1220 ( .A1(n1006), .A2(n1005), .Z(n1036) );
  or2 U1221 ( .A1(n431), .A2(n1307), .Z(n1462) );
  or2f U1222 ( .A1(n1032), .A2(n1081), .Z(n1002) );
  and2f U1223 ( .A1(n1446), .A2(n1032), .Z(n1034) );
  and2f U1224 ( .A1(n1437), .A2(n1469), .Z(n648) );
  or2f U1226 ( .A1(n1401), .A2(n1372), .Z(n1463) );
  or2f U1227 ( .A1(n1463), .A2(n1464), .Z(n76) );
  or2f U1228 ( .A1(n78), .A2(n141), .Z(n1464) );
  or2f U1229 ( .A1(n197), .A2(n1465), .Z(n172) );
  or2f U1230 ( .A1(n198), .A2(n862), .Z(n1465) );
  or2 U1231 ( .A1(n964), .A2(n1240), .Z(n914) );
  or2 U1232 ( .A1(n722), .A2(n159), .Z(n973) );
  and2f U1233 ( .A1(n1216), .A2(n989), .Z(n1466) );
  inv1f U1234 ( .I(n1466), .ZN(n1258) );
  inv1 U1235 ( .I(n989), .ZN(n1235) );
  inv1 U1236 ( .I(n1459), .ZN(n1230) );
  or2f U1237 ( .A1(n1005), .A2(q0), .Z(n976) );
  or2f U1238 ( .A1(n199), .A2(n200), .Z(n198) );
  or2 U1239 ( .A1(n1078), .A2(r0), .Z(n1287) );
  or2f U1240 ( .A1(n951), .A2(n802), .Z(n1078) );
  or2 U1241 ( .A1(n1133), .A2(n1441), .Z(n999) );
  and2 U1242 ( .A1(a0), .A2(r), .Z(n1468) );
  or2 U1243 ( .A1(n187), .A2(n796), .Z(n793) );
  and2f U1244 ( .A1(n317), .A2(n1067), .Z(n1404) );
  or2 U1246 ( .A1(n1451), .A2(n131), .Z(n1279) );
  and2f U1247 ( .A1(n1472), .A2(t), .Z(n1471) );
  inv1 U1248 ( .I(t), .ZN(n1210) );
  and2 U1249 ( .A1(w), .A2(n1235), .Z(n1237) );
  and2 U1250 ( .A1(y), .A2(n1235), .Z(n990) );
  and2 U1252 ( .A1(a), .A2(n421), .Z(n854) );
  and2 U1253 ( .A1(n284), .A2(n421), .Z(n1012) );
  and2 U1254 ( .A1(n616), .A2(n1258), .Z(n1259) );
  inv1 U1255 ( .I(n1032), .ZN(n1067) );
  and2 U1256 ( .A1(n1204), .A2(n1067), .Z(n473) );
  or2 U1257 ( .A1(n62), .A2(n1327), .Z(n1473) );
  or2f U1258 ( .A1(n1473), .A2(n1474), .Z(n1331) );
  or2 U1259 ( .A1(n1330), .A2(n133), .Z(n1474) );
  or2f U1260 ( .A1(n632), .A2(n1409), .Z(n1477) );
  or2 U1261 ( .A1(n1315), .A2(n1391), .Z(n1180) );
  or2f U1262 ( .A1(n1079), .A2(n960), .Z(n1133) );
  or2 U1263 ( .A1(n784), .A2(n785), .Z(n1478) );
  and2f U1264 ( .A1(e0), .A2(n1480), .Z(n1479) );
  inv1f U1265 ( .I(n1479), .ZN(n1079) );
  inv1f U1267 ( .I(u), .ZN(n1480) );
  or2 U1268 ( .A1(n1173), .A2(n174), .Z(n185) );
  or2f U1269 ( .A1(n1071), .A2(d0), .Z(n1491) );
  or2f U1270 ( .A1(n1470), .A2(n1491), .Z(n989) );
  or2 U1271 ( .A1(n1079), .A2(n1210), .Z(n1080) );
  or2 U1272 ( .A1(n77), .A2(n167), .Z(n163) );
  or2 U1273 ( .A1(n1333), .A2(n45), .Z(n1265) );
  or2f U1274 ( .A1(v), .A2(n1482), .Z(n1481) );
  inv1f U1275 ( .I(s), .ZN(n1482) );
  or2 U1276 ( .A1(n533), .A2(n534), .Z(n532) );
  and2 U1277 ( .A1(l), .A2(n317), .Z(n1095) );
  or2f U1278 ( .A1(n1495), .A2(n960), .Z(n1048) );
  or2f U1280 ( .A1(n1155), .A2(n1483), .Z(n1156) );
  and2 U1281 ( .A1(n1485), .A2(n1162), .Z(n1484) );
  or2 U1283 ( .A1(n1156), .A2(h0), .Z(n1186) );
  or2f U1284 ( .A1(n1166), .A2(m0), .Z(n916) );
  or2 U1285 ( .A1(n1156), .A2(n1487), .Z(n1301) );
  or2 U1286 ( .A1(h0), .A2(n870), .Z(n1487) );
  or2f U1287 ( .A1(n1156), .A2(n1493), .Z(n1492) );
  or2 U1288 ( .A1(n99), .A2(n367), .Z(n507) );
  or2 U1291 ( .A1(n119), .A2(n120), .Z(n118) );
  and2f U1292 ( .A1(n1390), .A2(n539), .Z(n564) );
  or2 U1293 ( .A1(n160), .A2(n131), .Z(n1488) );
  or2 U1296 ( .A1(h0), .A2(n1160), .Z(n1493) );
  or2f U1297 ( .A1(n1494), .A2(n1497), .Z(n1496) );
  inv1f U1298 ( .I(n1163), .ZN(n1497) );
  or2 U1299 ( .A1(n1327), .A2(n968), .Z(n1498) );
  or2f U1302 ( .A1(n916), .A2(n915), .Z(n1499) );
  or2f U1305 ( .A1(n1499), .A2(n1500), .Z(n951) );
  or2 U1306 ( .A1(n917), .A2(p0), .Z(n1500) );
  or2 U1307 ( .A1(n951), .A2(n931), .Z(n932) );
  inv1 U1311 ( .I(n1005), .ZN(n933) );
  or2 U1313 ( .A1(n1393), .A2(n1325), .Z(n1501) );
  inv1 U1314 ( .I(n0), .ZN(n1004) );
  and2 U1315 ( .A1(n1126), .A2(n1452), .Z(n657) );
  inv1 U1316 ( .I(n988), .ZN(n1366) );
  inv1 U1317 ( .I(n803), .ZN(n917) );
  and2 U1318 ( .A1(n1388), .A2(n1004), .Z(n803) );
  and2 U1319 ( .A1(n626), .A2(n849), .Z(n843) );
  and2 U1320 ( .A1(n548), .A2(c0), .Z(n849) );
  and2 U1322 ( .A1(n1390), .A2(n550), .Z(n263) );
  or2 U1323 ( .A1(n1388), .A2(n1004), .Z(n1006) );
  or2 U1324 ( .A1(n1354), .A2(n148), .Z(n146) );
  inv1 U1325 ( .I(n1068), .ZN(n1377) );
  or2 U1326 ( .A1(n1137), .A2(n1136), .Z(n1268) );
  or2 U1327 ( .A1(n246), .A2(n123), .Z(n1137) );
  or2 U1328 ( .A1(n247), .A2(n159), .Z(n1136) );
  or2 U1329 ( .A1(n1363), .A2(n1018), .Z(n1031) );
  or2 U1330 ( .A1(n597), .A2(n1379), .Z(n1018) );
  and2 U1331 ( .A1(n250), .A2(n), .Z(n68) );
  and2 U1332 ( .A1(n843), .A2(e), .Z(n175) );
  inv1 U1333 ( .I(n626), .ZN(n918) );
  inv1 U1336 ( .I(n966), .ZN(n1141) );
  or2 U1337 ( .A1(n965), .A2(n1019), .Z(n966) );
  or2 U1338 ( .A1(n1068), .A2(n1495), .Z(n965) );
  and2 U1339 ( .A1(n719), .A2(n1386), .Z(n716) );
  or2 U1341 ( .A1(n869), .A2(n1385), .Z(n373) );
  or2 U1342 ( .A1(n209), .A2(n210), .Z(n208) );
  or2 U1343 ( .A1(n1385), .A2(n1369), .Z(n210) );
  inv1 U1344 ( .I(n1070), .ZN(n1355) );
  or2 U1345 ( .A1(n1069), .A2(n1071), .Z(n1070) );
  or2 U1346 ( .A1(n1182), .A2(n1154), .Z(n1069) );
  or2 U1348 ( .A1(a0), .A2(n284), .Z(n338) );
  inv1 U1349 ( .I(c), .ZN(n325) );
  and2 U1350 ( .A1(z), .A2(l), .Z(n517) );
  or2 U1351 ( .A1(s0), .A2(o0), .Z(n802) );
  and2 U1352 ( .A1(x), .A2(f0), .Z(n1167) );
  and2 U1353 ( .A1(n1178), .A2(l0), .Z(n1157) );
  and2 U1354 ( .A1(n525), .A2(n899), .Z(n1083) );
  or2 U1355 ( .A1(d0), .A2(t), .Z(n947) );
  inv1 U1356 ( .I(n928), .ZN(n221) );
  or2 U1357 ( .A1(n1453), .A2(n1024), .Z(n928) );
  and2 U1358 ( .A1(n1434), .A2(n524), .Z(n872) );
  and2 U1359 ( .A1(e0), .A2(n525), .Z(n524) );
  inv1 U1361 ( .I(o), .ZN(n565) );
  and2 U1363 ( .A1(n1476), .A2(n1059), .Z(n1055) );
  and2 U1364 ( .A1(n1110), .A2(n1109), .Z(n1111) );
  and2 U1365 ( .A1(n1142), .A2(n1117), .Z(n1109) );
  and2 U1366 ( .A1(n1391), .A2(n1210), .Z(n1113) );
  and2 U1367 ( .A1(n1102), .A2(n1101), .Z(n312) );
  and2 U1368 ( .A1(n1210), .A2(n1100), .Z(n1101) );
  and2 U1369 ( .A1(n1148), .A2(n1099), .Z(n1102) );
  or2 U1370 ( .A1(n1117), .A2(c), .Z(n1100) );
  or2 U1371 ( .A1(n1390), .A2(c0), .Z(n940) );
  and2 U1372 ( .A1(n355), .A2(n356), .Z(n56) );
  and2 U1373 ( .A1(n1431), .A2(n1374), .Z(n355) );
  and2 U1376 ( .A1(n1386), .A2(y), .Z(n356) );
  inv1 U1378 ( .I(l), .ZN(n1392) );
  inv1 U1379 ( .I(n939), .ZN(n1372) );
  or2 U1381 ( .A1(n938), .A2(n937), .Z(n939) );
  or2 U1382 ( .A1(n936), .A2(n935), .Z(n937) );
  and2 U1386 ( .A1(n1083), .A2(n1374), .Z(n368) );
  inv1 U1387 ( .I(n1025), .ZN(n1360) );
  or2 U1388 ( .A1(n1024), .A2(n1023), .Z(n1025) );
  inv1 U1389 ( .I(n1476), .ZN(n1182) );
  or2 U1393 ( .A1(n1191), .A2(n1190), .Z(n1288) );
  or2 U1396 ( .A1(n999), .A2(n998), .Z(n1192) );
  or2 U1399 ( .A1(n997), .A2(n343), .Z(n998) );
  inv1 U1400 ( .I(n656), .ZN(n997) );
  and2 U1401 ( .A1(y), .A2(n473), .Z(n112) );
  inv1 U1406 ( .I(r), .ZN(n609) );
  and2 U1409 ( .A1(n550), .A2(a0), .Z(n790) );
  or2 U1410 ( .A1(n1355), .A2(n103), .Z(n97) );
  or2 U1415 ( .A1(n1366), .A2(n105), .Z(n103) );
  or2 U1416 ( .A1(n872), .A2(n221), .Z(n1267) );
  inv1 U1417 ( .I(n929), .ZN(n1375) );
  inv1 U1418 ( .I(n1275), .ZN(n1319) );
  or2 U1420 ( .A1(r), .A2(n1126), .Z(n1131) );
  and2 U1421 ( .A1(n424), .A2(n425), .Z(n862) );
  and2 U1424 ( .A1(n294), .A2(c), .Z(n424) );
  and2 U1425 ( .A1(n1442), .A2(n1238), .Z(n1243) );
  and2 U1427 ( .A1(a0), .A2(l), .Z(n616) );
  and2 U1428 ( .A1(n736), .A2(n696), .Z(n728) );
  and2 U1429 ( .A1(c0), .A2(n278), .Z(n736) );
  and2 U1434 ( .A1(n843), .A2(n844), .Z(n582) );
  and2 U1435 ( .A1(n279), .A2(n1431), .Z(n844) );
  inv1 U1436 ( .I(n1039), .ZN(n581) );
  or2 U1437 ( .A1(n1040), .A2(n1201), .Z(n1039) );
  or2 U1438 ( .A1(n871), .A2(n123), .Z(n624) );
  inv1 U1439 ( .I(n1082), .ZN(n223) );
  or2 U1440 ( .A1(n1217), .A2(n1081), .Z(n1082) );
  or2 U1442 ( .A1(n64), .A2(n216), .Z(n1307) );
  or2 U1443 ( .A1(n492), .A2(n1302), .Z(n1303) );
  and2 U1447 ( .A1(n493), .A2(n494), .Z(n492) );
  or2 U1448 ( .A1(n495), .A2(n496), .Z(n493) );
  and2 U1449 ( .A1(q), .A2(i), .Z(n496) );
  or2 U1450 ( .A1(n862), .A2(n1141), .Z(n230) );
  or2 U1451 ( .A1(n175), .A2(n591), .Z(n632) );
  and2 U1452 ( .A1(f), .A2(n389), .Z(n176) );
  and2 U1455 ( .A1(n390), .A2(n1376), .Z(n389) );
  inv1 U1456 ( .I(n1087), .ZN(n1352) );
  or2 U1457 ( .A1(n1086), .A2(n1214), .Z(n1087) );
  or2 U1460 ( .A1(n1315), .A2(a), .Z(n1086) );
  and2 U1461 ( .A1(n867), .A2(n1084), .Z(n866) );
  and2 U1462 ( .A1(n1431), .A2(y), .Z(n1084) );
  inv1 U1463 ( .I(n1085), .ZN(n867) );
  or2 U1464 ( .A1(n56), .A2(n866), .Z(n1412) );
  or2 U1466 ( .A1(n56), .A2(n57), .Z(n1410) );
  or2 U1467 ( .A1(n58), .A2(n59), .Z(n57) );
  or2 U1468 ( .A1(n871), .A2(n203), .Z(n1407) );
  or2 U1469 ( .A1(n528), .A2(n1362), .Z(n1037) );
  inv1 U1470 ( .I(n1192), .ZN(n1363) );
  and2 U1473 ( .A1(n476), .A2(n950), .Z(n777) );
  inv1 U1474 ( .I(r0), .ZN(n476) );
  and2 U1475 ( .A1(b0), .A2(n630), .Z(n123) );
  and2 U1476 ( .A1(n294), .A2(n631), .Z(n630) );
  or2 U1477 ( .A1(n209), .A2(n587), .Z(n165) );
  or2 U1478 ( .A1(n1325), .A2(n1403), .Z(n587) );
  or2 U1479 ( .A1(n68), .A2(n105), .Z(n249) );
  or2 U1480 ( .A1(n368), .A2(n369), .Z(n234) );
  or2 U1481 ( .A1(n223), .A2(n370), .Z(n369) );
  inv1 U1482 ( .I(n1285), .ZN(n370) );
  or2 U1487 ( .A1(n189), .A2(n190), .Z(n145) );
  or2 U1488 ( .A1(n1351), .A2(n191), .Z(n190) );
  or2 U1489 ( .A1(n192), .A2(n193), .Z(n189) );
  or2 U1490 ( .A1(n187), .A2(n188), .Z(n138) );
  or2 U1491 ( .A1(n1319), .A2(n182), .Z(n188) );
  and2 U1492 ( .A1(n1391), .A2(n278), .Z(n697) );
  inv1 U1493 ( .I(n1017), .ZN(n1379) );
  or2 U1494 ( .A1(n923), .A2(n922), .Z(n1017) );
  inv1 U1495 ( .I(p0), .ZN(n922) );
  or2 U1496 ( .A1(n1351), .A2(n168), .Z(n167) );
  or2 U1497 ( .A1(n112), .A2(n181), .Z(n177) );
  or2 U1498 ( .A1(n182), .A2(n1350), .Z(n181) );
  or2 U1499 ( .A1(n141), .A2(n142), .Z(n140) );
  or2 U1500 ( .A1(n157), .A2(n158), .Z(n154) );
  or2 U1501 ( .A1(n159), .A2(n160), .Z(n158) );
  inv1 U1502 ( .I(n1184), .ZN(n131) );
  or2 U1503 ( .A1(n1219), .A2(n1231), .Z(n1184) );
  or2 U1504 ( .A1(n1359), .A2(n1366), .Z(n132) );
  or2 U1505 ( .A1(n121), .A2(n122), .Z(n117) );
  or2 U1506 ( .A1(n123), .A2(n124), .Z(n122) );
  or2 U1507 ( .A1(n1189), .A2(n127), .Z(n126) );
  inv1 U1508 ( .I(n1188), .ZN(n1189) );
  or2 U1509 ( .A1(n1187), .A2(n1186), .Z(n1188) );
  and2 U1510 ( .A1(n1185), .A2(n1389), .Z(n1187) );
  and2 U1511 ( .A1(n1192), .A2(n1288), .Z(n1193) );
  or2 U1512 ( .A1(n1194), .A2(n1268), .Z(n1195) );
  or2 U1513 ( .A1(n112), .A2(n113), .Z(n108) );
  or2 U1514 ( .A1(n1359), .A2(n1350), .Z(n113) );
  inv1 U1515 ( .I(n1276), .ZN(n91) );
  or2 U1516 ( .A1(n1207), .A2(n1206), .Z(n64) );
  and2 U1517 ( .A1(n1458), .A2(n1205), .Z(n1206) );
  inv1 U1518 ( .I(n1203), .ZN(n1207) );
  and2 U1519 ( .A1(a0), .A2(n1204), .Z(n1205) );
  or2 U1520 ( .A1(n1319), .A2(n68), .Z(n1229) );
  or2 U1521 ( .A1(n1409), .A2(n1407), .Z(n50) );
  or2 U1522 ( .A1(n1261), .A2(n1255), .Z(n1398) );
  or2 U1523 ( .A1(n561), .A2(n175), .Z(n848) );
  inv1 U1524 ( .I(n903), .ZN(n1385) );
  or2 U1525 ( .A1(n902), .A2(n1495), .Z(n903) );
  and2 U1526 ( .A1(n1390), .A2(n525), .Z(n810) );
  inv1 U1527 ( .I(n906), .ZN(n1383) );
  or2 U1528 ( .A1(n905), .A2(n904), .Z(n906) );
  or2 U1529 ( .A1(n1096), .A2(n960), .Z(n905) );
  and2 U1530 ( .A1(n981), .A2(n1452), .Z(n982) );
  inv1 U1531 ( .I(n980), .ZN(n981) );
  or2 U1532 ( .A1(n1232), .A2(n1398), .Z(n808) );
  and2 U1533 ( .A1(n294), .A2(a), .Z(n1043) );
  inv1 U1534 ( .I(n1044), .ZN(n874) );
  or2 U1535 ( .A1(n575), .A2(n576), .Z(n1399) );
  or2 U1536 ( .A1(n1358), .A2(n578), .Z(n576) );
  or2 U1537 ( .A1(n579), .A2(n580), .Z(n575) );
  or2 U1538 ( .A1(n581), .A2(n582), .Z(n580) );
  or2 U1539 ( .A1(n572), .A2(n573), .Z(n571) );
  or2 U1540 ( .A1(n1141), .A2(n967), .Z(n968) );
  inv1 U1541 ( .I(n974), .ZN(n967) );
  inv1 U1542 ( .I(n1114), .ZN(n1380) );
  and2 U1543 ( .A1(n1472), .A2(e0), .Z(n1122) );
  and2 U1544 ( .A1(n1119), .A2(n1118), .Z(n1120) );
  or2 U1545 ( .A1(n1412), .A2(n1352), .Z(n348) );
  and2 U1546 ( .A1(n1361), .A2(n360), .Z(n347) );
  and2 U1547 ( .A1(n346), .A2(n343), .Z(n360) );
  or2 U1548 ( .A1(n875), .A2(n384), .Z(n214) );
  or2 U1549 ( .A1(n176), .A2(n1353), .Z(n384) );
  or2 U1550 ( .A1(n1147), .A2(n1146), .Z(n216) );
  and2 U1551 ( .A1(f), .A2(n1145), .Z(n1146) );
  and2 U1552 ( .A1(n483), .A2(n1211), .Z(n1147) );
  or2 U1553 ( .A1(n1370), .A2(n451), .Z(n483) );
  inv1 U1554 ( .I(n1106), .ZN(n900) );
  or2 U1555 ( .A1(n1350), .A2(n133), .Z(n1393) );
  and2 U1556 ( .A1(n278), .A2(n279), .Z(n277) );
  inv1 U1557 ( .I(k0), .ZN(n1178) );
  or2 U1558 ( .A1(n1059), .A2(n548), .Z(n957) );
  and2 U1559 ( .A1(n1210), .A2(n1148), .Z(n959) );
  or2 U1560 ( .A1(j0), .A2(i0), .Z(n870) );
  or2 U1561 ( .A1(n1104), .A2(n290), .Z(n289) );
  and2 U1562 ( .A1(a0), .A2(s), .Z(n290) );
  and2 U1563 ( .A1(x), .A2(n1108), .Z(n1104) );
  and2 U1564 ( .A1(n294), .A2(n1108), .Z(n1110) );
  and2 U1565 ( .A1(n281), .A2(s), .Z(n1107) );
  and2 U1566 ( .A1(n276), .A2(n277), .Z(n271) );
  and2 U1567 ( .A1(n1106), .A2(n1105), .Z(n272) );
  and2 U1568 ( .A1(c0), .A2(s), .Z(n276) );
  and2 U1569 ( .A1(n1210), .A2(n1088), .Z(n1094) );
  and2 U1570 ( .A1(n338), .A2(n1108), .Z(n1088) );
  and2 U1571 ( .A1(n323), .A2(n294), .Z(n1099) );
  or2 U1572 ( .A1(u), .A2(n325), .Z(n323) );
  inv1 U1573 ( .I(n1009), .ZN(n605) );
  or2 U1574 ( .A1(n1008), .A2(n1081), .Z(n1009) );
  inv1 U1575 ( .I(n1446), .ZN(n1001) );
  or2 U1576 ( .A1(y), .A2(n1081), .Z(n649) );
  or2 U1577 ( .A1(n652), .A2(w), .Z(n651) );
  inv1 U1578 ( .I(q0), .ZN(n1388) );
  inv1 U1579 ( .I(m0), .ZN(n935) );
  and2 U1580 ( .A1(n525), .A2(n1059), .Z(n1063) );
  inv1 U1581 ( .I(n1021), .ZN(n1064) );
  or2 U1582 ( .A1(n1020), .A2(n1019), .Z(n1021) );
  or2 U1583 ( .A1(n1441), .A2(n1495), .Z(n1020) );
  inv1 U1584 ( .I(n1083), .ZN(n1024) );
  and2 U1585 ( .A1(n1391), .A2(n548), .Z(n419) );
  or2 U1586 ( .A1(n151), .A2(n105), .Z(n150) );
  and2 U1587 ( .A1(n1391), .A2(x), .Z(n656) );
  inv1 U1588 ( .I(g0), .ZN(n1162) );
  or2 U1589 ( .A1(i0), .A2(n1185), .Z(n1160) );
  and2 U1590 ( .A1(n1285), .A2(n1284), .Z(n1286) );
  inv1 U1591 ( .I(n368), .ZN(n1284) );
  and2 U1592 ( .A1(n1289), .A2(n1288), .Z(n1290) );
  inv1 U1593 ( .I(n112), .ZN(n1289) );
  or2 U1594 ( .A1(n127), .A2(n1354), .Z(n243) );
  and2 U1595 ( .A1(z), .A2(n1392), .Z(n652) );
  inv1 U1596 ( .I(h0), .ZN(n1190) );
  inv1 U1597 ( .I(n947), .ZN(n948) );
  or2 U1598 ( .A1(n868), .A2(n1022), .Z(n1029) );
  and2 U1599 ( .A1(a0), .A2(n1064), .Z(n1022) );
  inv1 U1600 ( .I(k), .ZN(n1226) );
  inv1 U1601 ( .I(n1245), .ZN(n1238) );
  and2 U1602 ( .A1(n1392), .A2(n1126), .Z(n907) );
  and2 U1603 ( .A1(n317), .A2(a), .Z(n910) );
  and2 U1604 ( .A1(n732), .A2(c), .Z(n971) );
  and2 U1605 ( .A1(n294), .A2(a), .Z(n732) );
  inv1 U1606 ( .I(n832), .ZN(n913) );
  and2 U1607 ( .A1(n294), .A2(n325), .Z(n832) );
  inv1 U1608 ( .I(e), .ZN(n279) );
  or2 U1609 ( .A1(n963), .A2(n962), .Z(n753) );
  and2 U1610 ( .A1(n959), .A2(n958), .Z(n963) );
  and2 U1611 ( .A1(n1384), .A2(n1368), .Z(n962) );
  and2 U1612 ( .A1(n1472), .A2(n957), .Z(n958) );
  inv1 U1613 ( .I(q), .ZN(n497) );
  inv1 U1614 ( .I(n1158), .ZN(n1356) );
  inv1 U1615 ( .I(n961), .ZN(n1368) );
  or2 U1616 ( .A1(n960), .A2(n986), .Z(n961) );
  and2 U1617 ( .A1(n1210), .A2(n1374), .Z(n1053) );
  and2 U1618 ( .A1(n1142), .A2(n995), .Z(n674) );
  and2 U1619 ( .A1(n390), .A2(a), .Z(n995) );
  and2 U1620 ( .A1(n899), .A2(n1374), .Z(n1335) );
  and2 U1621 ( .A1(a0), .A2(t), .Z(n1336) );
  and2 U1622 ( .A1(n709), .A2(n1458), .Z(n1317) );
  inv1 U1623 ( .I(g), .ZN(n709) );
  and2 U1624 ( .A1(h), .A2(n497), .Z(n495) );
  and2 U1625 ( .A1(d), .A2(b0), .Z(n296) );
  inv1 U1626 ( .I(u), .ZN(n1117) );
  inv1 U1627 ( .I(n1008), .ZN(n1059) );
  and2 U1628 ( .A1(y), .A2(n1371), .Z(n58) );
  and2 U1629 ( .A1(n1374), .A2(a), .Z(n719) );
  inv1 U1630 ( .I(n854), .ZN(n996) );
  and2 U1631 ( .A1(n1067), .A2(n723), .Z(n871) );
  and2 U1632 ( .A1(a), .A2(n1367), .Z(n723) );
  and2 U1633 ( .A1(n1004), .A2(q0), .Z(n934) );
  inv1 U1634 ( .I(s0), .ZN(n931) );
  inv1 U1635 ( .I(o0), .ZN(n950) );
  inv1 U1636 ( .I(n1287), .ZN(n375) );
  and2 U1637 ( .A1(n1367), .A2(n1386), .Z(n105) );
  or2 U1638 ( .A1(n1360), .A2(n869), .Z(n1028) );
  or2 U1639 ( .A1(n1217), .A2(n1231), .Z(n1285) );
  and2 U1640 ( .A1(o), .A2(n410), .Z(n191) );
  and2 U1641 ( .A1(n1390), .A2(n1357), .Z(n410) );
  and2 U1642 ( .A1(n1168), .A2(n1167), .Z(n1169) );
  inv1 U1643 ( .I(b0), .ZN(n278) );
  and2 U1644 ( .A1(n420), .A2(n419), .Z(n1351) );
  and2 U1645 ( .A1(b0), .A2(n421), .Z(n420) );
  inv1 U1646 ( .I(a0), .ZN(n1081) );
  and2 U1647 ( .A1(n626), .A2(n419), .Z(n141) );
  inv1 U1648 ( .I(n1177), .ZN(n160) );
  or2 U1649 ( .A1(n1217), .A2(n1201), .Z(n1177) );
  or2 U1650 ( .A1(n1226), .A2(n451), .Z(n1231) );
  inv1 U1651 ( .I(j0), .ZN(n1185) );
  inv1 U1652 ( .I(i0), .ZN(n1389) );
  inv1 U1653 ( .I(n1011), .ZN(n1325) );
  or2 U1654 ( .A1(n1010), .A2(j), .Z(n1011) );
  or2 U1655 ( .A1(n1315), .A2(n1453), .Z(n1010) );
  inv1 U1656 ( .I(n930), .ZN(n85) );
  or2 U1657 ( .A1(n1153), .A2(n1315), .Z(n1275) );
  or2 U1658 ( .A1(n1441), .A2(n1154), .Z(n1153) );
  inv1 U1659 ( .I(n945), .ZN(n1369) );
  or2 U1660 ( .A1(n944), .A2(n947), .Z(n945) );
  or2 U1661 ( .A1(n943), .A2(n1198), .Z(n944) );
  or2 U1662 ( .A1(n1008), .A2(n1391), .Z(n943) );
  inv1 U1663 ( .I(n1073), .ZN(n1354) );
  or2 U1664 ( .A1(n1072), .A2(n1071), .Z(n1073) );
  or2 U1665 ( .A1(n1182), .A2(n1201), .Z(n1072) );
  or2 U1666 ( .A1(n1075), .A2(k), .Z(n1276) );
  or2 U1667 ( .A1(n1074), .A2(n451), .Z(n1075) );
  or2 U1668 ( .A1(n127), .A2(n105), .Z(n402) );
  or2 U1669 ( .A1(n1202), .A2(n1201), .Z(n1203) );
  and2 U1670 ( .A1(n1219), .A2(n1200), .Z(n1202) );
  or2 U1671 ( .A1(n1199), .A2(n1198), .Z(n1200) );
  inv1 U1672 ( .I(n1134), .ZN(n192) );
  or2 U1673 ( .A1(n1175), .A2(n1133), .Z(n1134) );
  and2 U1674 ( .A1(x), .A2(n1204), .Z(n1125) );
  and2 U1675 ( .A1(n910), .A2(n1129), .Z(n1261) );
  and2 U1676 ( .A1(v), .A2(n564), .Z(n250) );
  inv1 U1677 ( .I(d), .ZN(n294) );
  and2 U1678 ( .A1(n390), .A2(n842), .Z(n579) );
  and2 U1679 ( .A1(n664), .A2(n665), .Z(n578) );
  and2 U1680 ( .A1(a), .A2(n607), .Z(n665) );
  inv1 U1681 ( .I(n556), .ZN(n551) );
  and2 U1682 ( .A1(n557), .A2(n558), .Z(n556) );
  or2 U1683 ( .A1(h), .A2(q), .Z(n557) );
  or2 U1684 ( .A1(n497), .A2(i), .Z(n558) );
  or2 U1685 ( .A1(n552), .A2(n553), .Z(n494) );
  and2 U1686 ( .A1(n1054), .A2(n1053), .Z(n553) );
  and2 U1687 ( .A1(n1368), .A2(n1356), .Z(n552) );
  and2 U1688 ( .A1(c0), .A2(u), .Z(n1054) );
  and2 U1689 ( .A1(n1052), .A2(n1051), .Z(n559) );
  and2 U1690 ( .A1(p), .A2(n1142), .Z(n1052) );
  or2 U1691 ( .A1(n1050), .A2(n1145), .Z(n1051) );
  or2 U1692 ( .A1(n1397), .A2(n561), .Z(n560) );
  or2 U1693 ( .A1(n1058), .A2(n541), .Z(n540) );
  and2 U1694 ( .A1(n263), .A2(n), .Z(n541) );
  or2 U1695 ( .A1(n1339), .A2(n1338), .Z(n1340) );
  or2 U1696 ( .A1(n1337), .A2(n191), .Z(n1338) );
  or2 U1697 ( .A1(n1351), .A2(n1359), .Z(n1339) );
  and2 U1698 ( .A1(n1336), .A2(n1335), .Z(n1337) );
  or2 U1699 ( .A1(n200), .A2(n862), .Z(n1341) );
  inv1 U1700 ( .I(j), .ZN(n952) );
  or2 U1701 ( .A1(n1478), .A2(n511), .Z(n749) );
  or2 U1702 ( .A1(n45), .A2(n1379), .Z(n796) );
  or2 U1703 ( .A1(n1322), .A2(n1321), .Z(n1323) );
  and2 U1704 ( .A1(n1382), .A2(n970), .Z(n1322) );
  or2 U1705 ( .A1(n1320), .A2(n1319), .Z(n1321) );
  and2 U1706 ( .A1(n1318), .A2(n1317), .Z(n1320) );
  or2 U1707 ( .A1(n1326), .A2(n1360), .Z(n1330) );
  or2 U1708 ( .A1(n1325), .A2(n1387), .Z(n1326) );
  and2 U1709 ( .A1(n1113), .A2(n1112), .Z(n265) );
  and2 U1710 ( .A1(n296), .A2(n297), .Z(n260) );
  and2 U1711 ( .A1(n298), .A2(n1476), .Z(n297) );
  and2 U1712 ( .A1(u), .A2(n1471), .Z(n298) );
  or2 U1713 ( .A1(n920), .A2(n919), .Z(n1114) );
  or2 U1714 ( .A1(n918), .A2(c0), .Z(n919) );
  and2 U1715 ( .A1(n1117), .A2(n1432), .Z(n1118) );
  and2 U1716 ( .A1(n1391), .A2(n1116), .Z(n1119) );
  and2 U1717 ( .A1(n344), .A2(n343), .Z(n1116) );
  and2 U1718 ( .A1(t), .A2(n346), .Z(n344) );
  or2 U1719 ( .A1(n312), .A2(n313), .Z(n311) );
  or2 U1720 ( .A1(w), .A2(x), .Z(n346) );
  inv1 U1721 ( .I(b), .ZN(n343) );
  inv1 U1722 ( .I(z), .ZN(n451) );
  inv1 U1723 ( .I(n1246), .ZN(n1145) );
  or2 U1724 ( .A1(c0), .A2(n1142), .Z(n1106) );
  and2 U1725 ( .A1(n1151), .A2(n1458), .Z(n133) );
  and2 U1726 ( .A1(n1204), .A2(y), .Z(n1151) );
  or2 U1727 ( .A1(n1132), .A2(n1201), .Z(n1175) );
  and2 U1728 ( .A1(n1392), .A2(n1358), .Z(n1254) );
  and2 U1729 ( .A1(n609), .A2(e0), .Z(n608) );
  or2 U1730 ( .A1(n1278), .A2(n85), .Z(n1297) );
  inv1 U1731 ( .I(n1277), .ZN(n1278) );
  and2 U1732 ( .A1(n1276), .A2(n1275), .Z(n1277) );
  or2 U1733 ( .A1(n1272), .A2(n87), .Z(n1273) );
  or2 U1734 ( .A1(n1369), .A2(n81), .Z(n1272) );
  or2 U1735 ( .A1(n1269), .A2(n223), .Z(n1270) );
  or2 U1736 ( .A1(n1268), .A2(n142), .Z(n1269) );
  or2 U1737 ( .A1(n1375), .A2(n616), .Z(n638) );
  or2 U1738 ( .A1(n175), .A2(n176), .Z(n171) );
  and2 U1739 ( .A1(n250), .A2(n562), .Z(n1397) );
  inv1 U1740 ( .I(n563), .ZN(n562) );
  or2 U1741 ( .A1(n), .A2(m), .Z(n563) );
  or2 U1742 ( .A1(n1342), .A2(n65), .Z(n1343) );
  or2 U1743 ( .A1(n1341), .A2(n1340), .Z(n1342) );
  or2 U1744 ( .A1(n1304), .A2(n1303), .Z(n1309) );
  or2 U1745 ( .A1(n223), .A2(n1350), .Z(n1304) );
  or2 U1746 ( .A1(n229), .A2(n230), .Z(n225) );
  or2 U1747 ( .A1(n1359), .A2(n176), .Z(n229) );
  inv1 U1748 ( .I(n1248), .ZN(n1394) );
  or2 U1749 ( .A1(n1245), .A2(n1431), .Z(n1247) );
  inv1 U1750 ( .I(n1176), .ZN(n1350) );
  or2 U1751 ( .A1(n1175), .A2(n1489), .Z(n1176) );
  or2 U1752 ( .A1(n1410), .A2(n55), .Z(n51) );
  or2 U1753 ( .A1(n866), .A2(n1352), .Z(n52) );
  or2 U1754 ( .A1(n585), .A2(n586), .Z(n584) );
  or2 U1755 ( .A1(n119), .A2(n165), .Z(n586) );
  or2 U1756 ( .A1(n506), .A2(n507), .Z(e1) );
  or2 U1757 ( .A1(n123), .A2(n1363), .Z(n506) );
  or2 U1758 ( .A1(n121), .A2(n376), .Z(n361) );
  or2 U1759 ( .A1(n123), .A2(n242), .Z(n376) );
  or2 U1760 ( .A1(n148), .A2(n251), .Z(n232) );
  or2 U1761 ( .A1(n1355), .A2(n62), .Z(n251) );
  or2 U1762 ( .A1(n145), .A2(n138), .Z(n186) );
  or2 U1763 ( .A1(n177), .A2(n178), .Z(n161) );
  or2 U1764 ( .A1(n179), .A2(n1379), .Z(n178) );
  or2 U1765 ( .A1(n154), .A2(n155), .Z(n134) );
  or2 U1766 ( .A1(n1355), .A2(n156), .Z(n155) );
  or2 U1767 ( .A1(n115), .A2(n116), .Z(l1) );
  or2 U1768 ( .A1(n125), .A2(n126), .Z(n115) );
  or2 U1769 ( .A1(n131), .A2(n132), .Z(n125) );
  or2 U1770 ( .A1(n108), .A2(n109), .Z(n92) );
  inv1 U1771 ( .I(n1193), .ZN(n109) );
  or2 U1772 ( .A1(n62), .A2(n63), .Z(n61) );
  or2 U1773 ( .A1(n64), .A2(n65), .Z(n63) );
  or2 U1774 ( .A1(n45), .A2(n50), .Z(n1313) );
  or2 U1775 ( .A1(n1311), .A2(n1310), .Z(n1312) );
  or2 U1776 ( .A1(n1385), .A2(n591), .Z(n847) );
  or2 U1777 ( .A1(n1387), .A2(n848), .Z(n846) );
  or2 U1778 ( .A1(n808), .A2(n809), .Z(n725) );
  or2 U1779 ( .A1(n1383), .A2(n865), .Z(n809) );
  or2 U1780 ( .A1(n570), .A2(n571), .Z(n530) );
  or2 U1781 ( .A1(n1399), .A2(n873), .Z(n570) );
  or2 U1782 ( .A1(n347), .A2(n348), .Z(n252) );
  or2 U1783 ( .A1(n1387), .A2(n216), .Z(n215) );
  or2 U1784 ( .A1(n51), .A2(n52), .Z(t0) );
  or2 U1785 ( .A1(n861), .A2(n1358), .Z(a1) );
  or2 U1786 ( .A1(n1313), .A2(n1312), .Z(w1) );
  or2 U1787 ( .A1(n846), .A2(n847), .Z(a2) );
  or2 U1788 ( .A1(n252), .A2(n253), .Z(f2) );
  or2 U1789 ( .A1(n214), .A2(n215), .Z(h2) );
endmodule

