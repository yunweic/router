
module C1355_iscas ( o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, 
        a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, 
        d, c, b, a, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, 
        f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0 );
  input o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w,
         v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1,
         d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0;
  wire   n298, n299, n301, n302, n303, n304, n350, n386, n420, n463, n467,
         n476, n497, n498, n500, n501, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n520, n521, n522, n523, n524, n525,
         n526, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;

  and2 U283 ( .A1(n), .A2(n1021), .Z(n301) );
  and2 U287 ( .A1(p), .A2(n1019), .Z(n303) );
  and2 U336 ( .A1(l), .A2(n1018), .Z(n350) );
  and2 U381 ( .A1(i), .A2(n1021), .Z(n386) );
  and2 U422 ( .A1(j), .A2(n1020), .Z(n420) );
  and2 U476 ( .A1(k), .A2(n1019), .Z(n463) );
  and2 U507 ( .A1(k0), .A2(o0), .Z(n476) );
  or2 U524 ( .A1(n1017), .A2(n500), .Z(n498) );
  and2 U526 ( .A1(n500), .A2(n1017), .Z(n501) );
  and2 U540 ( .A1(n568), .A2(n508), .Z(n509) );
  inv1 U544 ( .I(k), .ZN(n512) );
  or2 U546 ( .A1(d0), .A2(n515), .Z(n514) );
  or2 U549 ( .A1(f0), .A2(n518), .Z(n517) );
  or2 U553 ( .A1(r), .A2(n522), .Z(n521) );
  or2 U555 ( .A1(s), .A2(n524), .Z(n523) );
  or2 U557 ( .A1(t), .A2(n526), .Z(n525) );
  or2 U560 ( .A1(n629), .A2(n628), .Z(n528) );
  or2 U562 ( .A1(q), .A2(n531), .Z(n530) );
  inv1 U564 ( .I(n1008), .ZN(n532) );
  inv1 U565 ( .I(n532), .ZN(n533) );
  or2 U566 ( .A1(c0), .A2(n535), .Z(n534) );
  inv1 U569 ( .I(n536), .ZN(n537) );
  or2 U570 ( .A1(e0), .A2(n539), .Z(n538) );
  inv1 U574 ( .I(y), .ZN(n974) );
  and2 U575 ( .A1(n974), .A2(u), .Z(n543) );
  and2 U577 ( .A1(y), .A2(n946), .Z(n542) );
  or2 U578 ( .A1(n543), .A2(n542), .Z(n500) );
  inv1 U579 ( .I(q), .ZN(n927) );
  and2 U580 ( .A1(n927), .A2(c0), .Z(n545) );
  inv1 U581 ( .I(c0), .ZN(n1001) );
  and2 U582 ( .A1(q), .A2(n1001), .Z(n544) );
  or2 U583 ( .A1(n545), .A2(n544), .Z(n546) );
  inv1 U584 ( .I(n546), .ZN(n1017) );
  inv1 U586 ( .I(o), .ZN(n1019) );
  inv1 U587 ( .I(n), .ZN(n1020) );
  inv1 U588 ( .I(m), .ZN(n1021) );
  inv1 U589 ( .I(p), .ZN(n1018) );
  and2 U591 ( .A1(n547), .A2(n476), .Z(n550) );
  inv1 U592 ( .I(n476), .ZN(n548) );
  or2 U594 ( .A1(n550), .A2(n549), .Z(n574) );
  or2 U599 ( .A1(n552), .A2(n551), .Z(n556) );
  inv1 U605 ( .I(n557), .ZN(n555) );
  and2 U606 ( .A1(n556), .A2(n555), .Z(n560) );
  inv1 U607 ( .I(n556), .ZN(n558) );
  and2 U612 ( .A1(n863), .A2(h), .Z(n562) );
  and2 U613 ( .A1(n516), .A2(g), .Z(n561) );
  inv1 U615 ( .I(e), .ZN(n853) );
  and2 U616 ( .A1(f), .A2(n853), .Z(n564) );
  inv1 U617 ( .I(f), .ZN(n858) );
  and2 U618 ( .A1(n858), .A2(e), .Z(n563) );
  or2 U619 ( .A1(n564), .A2(n563), .Z(n567) );
  inv1 U620 ( .I(n567), .ZN(n565) );
  inv1 U622 ( .I(n566), .ZN(n568) );
  and2 U623 ( .A1(n568), .A2(n508), .Z(n569) );
  and2 U625 ( .A1(n600), .A2(n510), .Z(n572) );
  inv1 U626 ( .I(n631), .ZN(n630) );
  or2 U628 ( .A1(n572), .A2(n571), .Z(n575) );
  inv1 U629 ( .I(n575), .ZN(n573) );
  and2 U630 ( .A1(n574), .A2(n573), .Z(n578) );
  inv1 U631 ( .I(n574), .ZN(n576) );
  inv1 U634 ( .I(a0), .ZN(n984) );
  and2 U635 ( .A1(n984), .A2(e0), .Z(n580) );
  inv1 U636 ( .I(e0), .ZN(n1009) );
  and2 U637 ( .A1(a0), .A2(n1009), .Z(n579) );
  or2 U638 ( .A1(n580), .A2(n579), .Z(n584) );
  inv1 U639 ( .I(s), .ZN(n933) );
  and2 U640 ( .A1(n933), .A2(w), .Z(n582) );
  inv1 U641 ( .I(w), .ZN(n956) );
  and2 U642 ( .A1(s), .A2(n956), .Z(n581) );
  or2 U643 ( .A1(n582), .A2(n581), .Z(n585) );
  inv1 U644 ( .I(n585), .ZN(n583) );
  and2 U645 ( .A1(n584), .A2(n583), .Z(n588) );
  inv1 U646 ( .I(n584), .ZN(n586) );
  and2 U647 ( .A1(n586), .A2(n585), .Z(n587) );
  or2 U648 ( .A1(n588), .A2(n587), .Z(n611) );
  inv1 U649 ( .I(o0), .ZN(n808) );
  inv1 U650 ( .I(m0), .ZN(n589) );
  or2 U651 ( .A1(n808), .A2(n589), .Z(n605) );
  and2 U653 ( .A1(k), .A2(n893), .Z(n591) );
  and2 U654 ( .A1(n512), .A2(l), .Z(n590) );
  or2 U655 ( .A1(n591), .A2(n590), .Z(n595) );
  inv1 U656 ( .I(i), .ZN(n878) );
  and2 U657 ( .A1(j), .A2(n878), .Z(n593) );
  and2 U666 ( .A1(n513), .A2(n600), .Z(n603) );
  inv1 U667 ( .I(n658), .ZN(n660) );
  and2 U668 ( .A1(n660), .A2(n601), .Z(n602) );
  and2 U671 ( .A1(n605), .A2(n604), .Z(n609) );
  inv1 U672 ( .I(n605), .ZN(n606) );
  and2 U673 ( .A1(n607), .A2(n606), .Z(n608) );
  inv1 U675 ( .I(n612), .ZN(n610) );
  inv1 U677 ( .I(n611), .ZN(n613) );
  inv1 U681 ( .I(b0), .ZN(n990) );
  and2 U682 ( .A1(n990), .A2(f0), .Z(n617) );
  inv1 U683 ( .I(f0), .ZN(n1014) );
  and2 U684 ( .A1(b0), .A2(n1014), .Z(n616) );
  or2 U685 ( .A1(n617), .A2(n616), .Z(n621) );
  and2 U687 ( .A1(n937), .A2(x), .Z(n619) );
  and2 U689 ( .A1(t), .A2(n962), .Z(n618) );
  or2 U690 ( .A1(n619), .A2(n618), .Z(n622) );
  inv1 U691 ( .I(n622), .ZN(n620) );
  and2 U692 ( .A1(n621), .A2(n620), .Z(n625) );
  inv1 U693 ( .I(n621), .ZN(n623) );
  and2 U694 ( .A1(n623), .A2(n622), .Z(n624) );
  or2 U695 ( .A1(n625), .A2(n624), .Z(n642) );
  inv1 U696 ( .I(n298), .ZN(n626) );
  and2 U697 ( .A1(n626), .A2(n299), .Z(n629) );
  inv1 U698 ( .I(n299), .ZN(n627) );
  inv1 U702 ( .I(n659), .ZN(n657) );
  and2 U703 ( .A1(n657), .A2(n510), .Z(n632) );
  inv1 U705 ( .I(n0), .ZN(n634) );
  or2 U706 ( .A1(n808), .A2(n634), .Z(n637) );
  inv1 U707 ( .I(n637), .ZN(n635) );
  inv1 U709 ( .I(n636), .ZN(n638) );
  inv1 U714 ( .I(n642), .ZN(n644) );
  and2 U715 ( .A1(n644), .A2(n643), .Z(n645) );
  or2 U718 ( .A1(n919), .A2(n540), .Z(n827) );
  inv1 U719 ( .I(z), .ZN(n979) );
  and2 U720 ( .A1(n979), .A2(d0), .Z(n648) );
  inv1 U721 ( .I(d0), .ZN(n1005) );
  and2 U722 ( .A1(z), .A2(n1005), .Z(n647) );
  or2 U723 ( .A1(n648), .A2(n647), .Z(n652) );
  and2 U725 ( .A1(n930), .A2(v), .Z(n650) );
  inv1 U726 ( .I(v), .ZN(n951) );
  and2 U727 ( .A1(r), .A2(n951), .Z(n649) );
  or2 U728 ( .A1(n650), .A2(n649), .Z(n653) );
  inv1 U729 ( .I(n653), .ZN(n651) );
  and2 U730 ( .A1(n652), .A2(n651), .Z(n656) );
  inv1 U731 ( .I(n652), .ZN(n654) );
  and2 U732 ( .A1(n654), .A2(n653), .Z(n655) );
  or2 U733 ( .A1(n656), .A2(n655), .Z(n671) );
  and2 U734 ( .A1(n513), .A2(n657), .Z(n662) );
  inv1 U737 ( .I(l0), .ZN(n663) );
  or2 U738 ( .A1(n808), .A2(n663), .Z(n666) );
  inv1 U739 ( .I(n666), .ZN(n664) );
  inv1 U746 ( .I(n671), .ZN(n673) );
  and2 U747 ( .A1(n673), .A2(n672), .Z(n674) );
  and2 U750 ( .A1(e), .A2(n829), .Z(n677) );
  and2 U751 ( .A1(n853), .A2(a), .Z(n676) );
  or2 U752 ( .A1(n677), .A2(n676), .Z(n688) );
  and2 U753 ( .A1(n956), .A2(x), .Z(n679) );
  and2 U754 ( .A1(w), .A2(n962), .Z(n678) );
  or2 U755 ( .A1(n679), .A2(n678), .Z(n683) );
  and2 U756 ( .A1(v), .A2(n946), .Z(n681) );
  inv1 U759 ( .I(n684), .ZN(n682) );
  and2 U760 ( .A1(n683), .A2(n682), .Z(n687) );
  inv1 U761 ( .I(n683), .ZN(n685) );
  and2 U765 ( .A1(n688), .A2(n776), .Z(n691) );
  inv1 U766 ( .I(n688), .ZN(n689) );
  and2 U767 ( .A1(n689), .A2(n774), .Z(n690) );
  or2 U768 ( .A1(n691), .A2(n690), .Z(n715) );
  or2 U771 ( .A1(n693), .A2(n692), .Z(n697) );
  inv1 U775 ( .I(n698), .ZN(n696) );
  and2 U776 ( .A1(n697), .A2(n696), .Z(n701) );
  inv1 U777 ( .I(n697), .ZN(n699) );
  and2 U780 ( .A1(n878), .A2(m), .Z(n702) );
  or2 U781 ( .A1(n702), .A2(n386), .Z(n704) );
  inv1 U782 ( .I(n704), .ZN(n703) );
  and2 U783 ( .A1(n738), .A2(n703), .Z(n706) );
  inv1 U784 ( .I(n738), .ZN(n740) );
  and2 U785 ( .A1(n740), .A2(n704), .Z(n705) );
  or2 U786 ( .A1(n706), .A2(n705), .Z(n709) );
  inv1 U787 ( .I(g0), .ZN(n707) );
  or2 U788 ( .A1(n707), .A2(n808), .Z(n710) );
  inv1 U789 ( .I(n710), .ZN(n708) );
  and2 U790 ( .A1(n709), .A2(n708), .Z(n713) );
  inv1 U791 ( .I(n709), .ZN(n711) );
  and2 U792 ( .A1(n711), .A2(n710), .Z(n712) );
  or2 U793 ( .A1(n713), .A2(n712), .Z(n716) );
  inv1 U794 ( .I(n716), .ZN(n714) );
  inv1 U796 ( .I(n715), .ZN(n717) );
  and2 U797 ( .A1(n717), .A2(n716), .Z(n718) );
  and2 U799 ( .A1(b0), .A2(n984), .Z(n721) );
  and2 U800 ( .A1(n990), .A2(a0), .Z(n720) );
  or2 U801 ( .A1(n721), .A2(n720), .Z(n725) );
  and2 U802 ( .A1(z), .A2(n974), .Z(n723) );
  and2 U803 ( .A1(n979), .A2(y), .Z(n722) );
  or2 U804 ( .A1(n723), .A2(n722), .Z(n726) );
  inv1 U805 ( .I(n726), .ZN(n724) );
  and2 U806 ( .A1(n725), .A2(n724), .Z(n729) );
  inv1 U807 ( .I(n725), .ZN(n727) );
  and2 U811 ( .A1(g), .A2(n839), .Z(n731) );
  and2 U812 ( .A1(n863), .A2(c), .Z(n730) );
  or2 U813 ( .A1(n731), .A2(n730), .Z(n732) );
  and2 U814 ( .A1(n804), .A2(n732), .Z(n735) );
  inv1 U815 ( .I(n732), .ZN(n733) );
  and2 U816 ( .A1(n802), .A2(n733), .Z(n734) );
  or2 U817 ( .A1(n735), .A2(n734), .Z(n751) );
  and2 U818 ( .A1(n512), .A2(o), .Z(n736) );
  or2 U819 ( .A1(n736), .A2(n463), .Z(n739) );
  inv1 U820 ( .I(n739), .ZN(n737) );
  and2 U821 ( .A1(n738), .A2(n737), .Z(n742) );
  and2 U822 ( .A1(n740), .A2(n739), .Z(n741) );
  or2 U823 ( .A1(n742), .A2(n741), .Z(n745) );
  inv1 U824 ( .I(i0), .ZN(n743) );
  or2 U825 ( .A1(n808), .A2(n743), .Z(n746) );
  inv1 U826 ( .I(n746), .ZN(n744) );
  and2 U827 ( .A1(n745), .A2(n744), .Z(n749) );
  inv1 U828 ( .I(n745), .ZN(n747) );
  and2 U829 ( .A1(n747), .A2(n746), .Z(n748) );
  or2 U830 ( .A1(n749), .A2(n748), .Z(n752) );
  inv1 U831 ( .I(n752), .ZN(n750) );
  inv1 U833 ( .I(n751), .ZN(n753) );
  and2 U834 ( .A1(n753), .A2(n752), .Z(n754) );
  and2 U837 ( .A1(f0), .A2(n1009), .Z(n757) );
  and2 U838 ( .A1(n1014), .A2(e0), .Z(n756) );
  or2 U839 ( .A1(n757), .A2(n756), .Z(n761) );
  and2 U840 ( .A1(d0), .A2(n1001), .Z(n759) );
  and2 U841 ( .A1(n1005), .A2(c0), .Z(n758) );
  or2 U842 ( .A1(n759), .A2(n758), .Z(n762) );
  inv1 U843 ( .I(n762), .ZN(n760) );
  and2 U844 ( .A1(n761), .A2(n760), .Z(n765) );
  inv1 U845 ( .I(n761), .ZN(n763) );
  and2 U846 ( .A1(n763), .A2(n762), .Z(n764) );
  or2 U847 ( .A1(n765), .A2(n764), .Z(n796) );
  inv1 U848 ( .I(n796), .ZN(n794) );
  and2 U849 ( .A1(h), .A2(n845), .Z(n767) );
  and2 U850 ( .A1(n516), .A2(d), .Z(n766) );
  or2 U851 ( .A1(n767), .A2(n766), .Z(n768) );
  and2 U852 ( .A1(n794), .A2(n768), .Z(n771) );
  inv1 U853 ( .I(n768), .ZN(n769) );
  and2 U854 ( .A1(n796), .A2(n769), .Z(n770) );
  or2 U855 ( .A1(n771), .A2(n770), .Z(n787) );
  and2 U856 ( .A1(n893), .A2(p), .Z(n772) );
  or2 U857 ( .A1(n772), .A2(n350), .Z(n775) );
  inv1 U858 ( .I(n775), .ZN(n773) );
  and2 U859 ( .A1(n774), .A2(n773), .Z(n778) );
  and2 U860 ( .A1(n776), .A2(n775), .Z(n777) );
  or2 U861 ( .A1(n778), .A2(n777), .Z(n781) );
  inv1 U862 ( .I(j0), .ZN(n779) );
  or2 U863 ( .A1(n808), .A2(n779), .Z(n782) );
  inv1 U864 ( .I(n782), .ZN(n780) );
  and2 U865 ( .A1(n781), .A2(n780), .Z(n785) );
  inv1 U866 ( .I(n781), .ZN(n783) );
  and2 U867 ( .A1(n783), .A2(n782), .Z(n784) );
  inv1 U869 ( .I(n788), .ZN(n786) );
  inv1 U871 ( .I(n787), .ZN(n789) );
  and2 U874 ( .A1(f), .A2(n834), .Z(n793) );
  and2 U875 ( .A1(n858), .A2(b), .Z(n792) );
  or2 U876 ( .A1(n793), .A2(n792), .Z(n795) );
  and2 U877 ( .A1(n795), .A2(n794), .Z(n799) );
  inv1 U878 ( .I(n795), .ZN(n797) );
  and2 U879 ( .A1(n797), .A2(n796), .Z(n798) );
  or2 U880 ( .A1(n799), .A2(n798), .Z(n816) );
  and2 U881 ( .A1(n883), .A2(n), .Z(n800) );
  or2 U882 ( .A1(n800), .A2(n420), .Z(n803) );
  inv1 U883 ( .I(n803), .ZN(n801) );
  and2 U885 ( .A1(n804), .A2(n803), .Z(n805) );
  or2 U886 ( .A1(n806), .A2(n805), .Z(n810) );
  inv1 U887 ( .I(h0), .ZN(n807) );
  or2 U888 ( .A1(n808), .A2(n807), .Z(n811) );
  inv1 U889 ( .I(n811), .ZN(n809) );
  and2 U890 ( .A1(n810), .A2(n809), .Z(n814) );
  and2 U892 ( .A1(n812), .A2(n811), .Z(n813) );
  inv1 U894 ( .I(n817), .ZN(n815) );
  inv1 U896 ( .I(n816), .ZN(n818) );
  inv1 U909 ( .I(n830), .ZN(n828) );
  or2 U910 ( .A1(n828), .A2(a), .Z(n832) );
  or2 U911 ( .A1(n830), .A2(n829), .Z(n831) );
  and2 U912 ( .A1(n832), .A2(n831), .Z(p0) );
  inv1 U914 ( .I(n835), .ZN(n833) );
  or2 U915 ( .A1(n833), .A2(b), .Z(n837) );
  and2 U917 ( .A1(n837), .A2(n836), .Z(q0) );
  inv1 U919 ( .I(n840), .ZN(n838) );
  or2 U920 ( .A1(n838), .A2(c), .Z(n842) );
  and2 U922 ( .A1(n842), .A2(n841), .Z(r0) );
  or2 U925 ( .A1(n844), .A2(d), .Z(n848) );
  or2 U926 ( .A1(n846), .A2(n845), .Z(n847) );
  and2 U927 ( .A1(n848), .A2(n847), .Z(s0) );
  or2 U929 ( .A1(n850), .A2(n536), .Z(n851) );
  or2 U934 ( .A1(n852), .A2(e), .Z(n856) );
  or2 U935 ( .A1(n854), .A2(n853), .Z(n855) );
  and2 U936 ( .A1(n856), .A2(n855), .Z(t0) );
  or2 U939 ( .A1(n857), .A2(f), .Z(n861) );
  or2 U940 ( .A1(n859), .A2(n858), .Z(n860) );
  and2 U941 ( .A1(n861), .A2(n860), .Z(u0) );
  or2 U944 ( .A1(n862), .A2(g), .Z(n866) );
  or2 U945 ( .A1(n864), .A2(n863), .Z(n865) );
  and2 U946 ( .A1(n866), .A2(n865), .Z(v0) );
  or2 U949 ( .A1(n868), .A2(h), .Z(n871) );
  or2 U950 ( .A1(n869), .A2(n516), .Z(n870) );
  and2 U951 ( .A1(n871), .A2(n870), .Z(w0) );
  inv1 U952 ( .I(n1000), .ZN(n897) );
  or2 U953 ( .A1(n533), .A2(n537), .Z(n872) );
  or2 U954 ( .A1(n897), .A2(n872), .Z(n876) );
  inv1 U958 ( .I(n879), .ZN(n877) );
  or2 U959 ( .A1(n877), .A2(i), .Z(n881) );
  or2 U960 ( .A1(n879), .A2(n878), .Z(n880) );
  and2 U961 ( .A1(n881), .A2(n880), .Z(x0) );
  inv1 U963 ( .I(n884), .ZN(n882) );
  or2 U964 ( .A1(n882), .A2(j), .Z(n886) );
  and2 U966 ( .A1(n886), .A2(n885), .Z(y0) );
  or2 U970 ( .A1(k), .A2(n888), .Z(n889) );
  and2 U971 ( .A1(n890), .A2(n889), .Z(z0) );
  or2 U974 ( .A1(n892), .A2(l), .Z(n896) );
  or2 U975 ( .A1(n894), .A2(n893), .Z(n895) );
  and2 U976 ( .A1(n896), .A2(n895), .Z(a1) );
  or2 U977 ( .A1(n917), .A2(n897), .Z(n899) );
  or2 U981 ( .A1(n900), .A2(m), .Z(n903) );
  or2 U982 ( .A1(n901), .A2(n1021), .Z(n902) );
  and2 U983 ( .A1(n903), .A2(n902), .Z(b1) );
  or2 U986 ( .A1(n904), .A2(n), .Z(n907) );
  or2 U987 ( .A1(n905), .A2(n1020), .Z(n906) );
  and2 U988 ( .A1(n907), .A2(n906), .Z(c1) );
  or2 U991 ( .A1(n908), .A2(o), .Z(n911) );
  or2 U992 ( .A1(n909), .A2(n1019), .Z(n910) );
  and2 U993 ( .A1(n911), .A2(n910), .Z(d1) );
  or2 U996 ( .A1(n913), .A2(p), .Z(n916) );
  or2 U997 ( .A1(n914), .A2(n1018), .Z(n915) );
  and2 U998 ( .A1(n916), .A2(n915), .Z(e1) );
  and2 U1000 ( .A1(n533), .A2(n918), .Z(n922) );
  and2 U1002 ( .A1(n537), .A2(n920), .Z(n921) );
  or2 U1008 ( .A1(n924), .A2(n1023), .Z(n925) );
  or2 U1011 ( .A1(n928), .A2(n927), .Z(n929) );
  and2 U1012 ( .A1(n530), .A2(n929), .Z(f1) );
  or2 U1014 ( .A1(n931), .A2(n930), .Z(n932) );
  and2 U1015 ( .A1(n521), .A2(n932), .Z(g1) );
  or2 U1017 ( .A1(n934), .A2(n933), .Z(n935) );
  and2 U1018 ( .A1(n523), .A2(n935), .Z(h1) );
  and2 U1021 ( .A1(n525), .A2(n939), .Z(i1) );
  inv1 U1022 ( .I(n969), .ZN(n994) );
  or2 U1023 ( .A1(n1025), .A2(n994), .Z(n941) );
  or2 U1025 ( .A1(n1028), .A2(n1024), .Z(n943) );
  or2 U1029 ( .A1(n945), .A2(u), .Z(n949) );
  or2 U1030 ( .A1(n947), .A2(n946), .Z(n948) );
  and2 U1031 ( .A1(n949), .A2(n948), .Z(j1) );
  or2 U1034 ( .A1(n950), .A2(v), .Z(n954) );
  or2 U1035 ( .A1(n952), .A2(n951), .Z(n953) );
  and2 U1036 ( .A1(n954), .A2(n953), .Z(k1) );
  or2 U1039 ( .A1(n955), .A2(w), .Z(n959) );
  or2 U1040 ( .A1(n957), .A2(n956), .Z(n958) );
  and2 U1041 ( .A1(n959), .A2(n958), .Z(l1) );
  or2 U1044 ( .A1(n961), .A2(x), .Z(n965) );
  or2 U1045 ( .A1(n963), .A2(n962), .Z(n964) );
  and2 U1046 ( .A1(n965), .A2(n964), .Z(m1) );
  or2 U1048 ( .A1(n1027), .A2(n1023), .Z(n968) );
  or2 U1050 ( .A1(n1026), .A2(n969), .Z(n971) );
  or2 U1054 ( .A1(n973), .A2(y), .Z(n977) );
  or2 U1055 ( .A1(n975), .A2(n974), .Z(n976) );
  and2 U1056 ( .A1(n977), .A2(n976), .Z(n1) );
  or2 U1059 ( .A1(n978), .A2(z), .Z(n982) );
  or2 U1060 ( .A1(n980), .A2(n979), .Z(n981) );
  and2 U1061 ( .A1(n982), .A2(n981), .Z(o1) );
  or2 U1064 ( .A1(n983), .A2(a0), .Z(n987) );
  or2 U1065 ( .A1(n985), .A2(n984), .Z(n986) );
  and2 U1066 ( .A1(n987), .A2(n986), .Z(p1) );
  or2 U1069 ( .A1(n989), .A2(b0), .Z(n993) );
  or2 U1070 ( .A1(n991), .A2(n990), .Z(n992) );
  and2 U1071 ( .A1(n993), .A2(n992), .Z(q1) );
  or2 U1073 ( .A1(n997), .A2(n1027), .Z(n998) );
  or2 U1076 ( .A1(n1002), .A2(n1001), .Z(n1003) );
  and2 U1077 ( .A1(n534), .A2(n1003), .Z(r1) );
  or2 U1079 ( .A1(n1006), .A2(n1005), .Z(n1007) );
  and2 U1080 ( .A1(n514), .A2(n1007), .Z(s1) );
  or2 U1082 ( .A1(n1010), .A2(n1009), .Z(n1011) );
  and2 U1083 ( .A1(n538), .A2(n1011), .Z(t1) );
  or2 U1085 ( .A1(n1015), .A2(n1014), .Z(n1016) );
  and2 U1086 ( .A1(n517), .A2(n1016), .Z(u1) );
  inv1f U538 ( .I(n854), .ZN(n852) );
  inv1f U539 ( .I(n859), .ZN(n857) );
  inv1f U541 ( .I(n901), .ZN(n900) );
  inv1f U542 ( .I(n905), .ZN(n904) );
  inv1f U543 ( .I(n869), .ZN(n868) );
  inv1f U545 ( .I(n914), .ZN(n913) );
  inv1f U547 ( .I(n864), .ZN(n862) );
  inv1f U548 ( .I(n909), .ZN(n908) );
  or2 U550 ( .A1(n876), .A2(n969), .Z(n1022) );
  inv1 U551 ( .I(n887), .ZN(n888) );
  or2 U552 ( .A1(n1022), .A2(n875), .Z(n887) );
  inv1f U554 ( .I(n963), .ZN(n961) );
  inv1f U556 ( .I(n991), .ZN(n989) );
  inv1f U558 ( .I(n957), .ZN(n955) );
  inv1f U559 ( .I(n985), .ZN(n983) );
  inv1f U561 ( .I(n952), .ZN(n950) );
  inv1f U563 ( .I(n980), .ZN(n978) );
  inv1f U567 ( .I(n947), .ZN(n945) );
  inv1f U568 ( .I(n975), .ZN(n973) );
  inv1f U571 ( .I(n938), .ZN(n526) );
  inv1f U572 ( .I(n1015), .ZN(n518) );
  inv1f U573 ( .I(n934), .ZN(n524) );
  inv1f U576 ( .I(n1010), .ZN(n539) );
  inv1f U585 ( .I(n931), .ZN(n522) );
  inv1f U590 ( .I(n1006), .ZN(n515) );
  inv1f U593 ( .I(n928), .ZN(n531) );
  inv1f U595 ( .I(n1002), .ZN(n535) );
  inv1 U596 ( .I(b), .ZN(n834) );
  inv1 U597 ( .I(j), .ZN(n883) );
  and2 U598 ( .A1(n883), .A2(i), .Z(n592) );
  and2 U600 ( .A1(n951), .A2(u), .Z(n680) );
  and2 U601 ( .A1(c), .A2(n845), .Z(n552) );
  and2 U602 ( .A1(n839), .A2(d), .Z(n551) );
  inv1 U603 ( .I(n802), .ZN(n804) );
  inv1 U604 ( .I(n601), .ZN(n600) );
  inv1 U608 ( .I(n467), .ZN(n547) );
  inv1 U609 ( .I(a), .ZN(n829) );
  inv1 U610 ( .I(d), .ZN(n845) );
  inv1 U611 ( .I(g), .ZN(n863) );
  inv1 U614 ( .I(l), .ZN(n893) );
  inv1 U621 ( .I(u), .ZN(n946) );
  inv1 U624 ( .I(x), .ZN(n962) );
  or2 U627 ( .A1(n835), .A2(n834), .Z(n836) );
  or2 U632 ( .A1(n840), .A2(n839), .Z(n841) );
  or2 U633 ( .A1(n884), .A2(n883), .Z(n885) );
  inv1f U652 ( .I(n774), .ZN(n776) );
  or2f U658 ( .A1(n942), .A2(n970), .Z(n997) );
  or2f U659 ( .A1(n791), .A2(n790), .Z(n942) );
  or2f U660 ( .A1(n1000), .A2(n1008), .Z(n919) );
  or2f U661 ( .A1(n615), .A2(n614), .Z(n1008) );
  inv1f U662 ( .I(c), .ZN(n839) );
  and2f U663 ( .A1(b), .A2(n829), .Z(n554) );
  and2f U664 ( .A1(n834), .A2(a), .Z(n553) );
  and2 U665 ( .A1(n802), .A2(n801), .Z(n806) );
  and2 U669 ( .A1(n497), .A2(n498), .Z(n467) );
  inv1 U670 ( .I(n501), .ZN(n497) );
  and2 U674 ( .A1(n576), .A2(n575), .Z(n577) );
  or2 U676 ( .A1(n593), .A2(n592), .Z(n596) );
  and2 U678 ( .A1(n1018), .A2(o), .Z(n304) );
  inv1 U679 ( .I(n810), .ZN(n812) );
  or2 U680 ( .A1(n687), .A2(n686), .Z(n774) );
  or2 U686 ( .A1(n562), .A2(n561), .Z(n566) );
  or2 U688 ( .A1(n603), .A2(n602), .Z(n607) );
  or2 U699 ( .A1(n554), .A2(n553), .Z(n557) );
  and2 U700 ( .A1(n727), .A2(n726), .Z(n728) );
  and2 U701 ( .A1(n715), .A2(n714), .Z(n719) );
  and2 U704 ( .A1(n787), .A2(n786), .Z(n791) );
  and2 U708 ( .A1(n789), .A2(n788), .Z(n790) );
  inv1 U710 ( .I(n672), .ZN(n670) );
  and2 U711 ( .A1(n467), .A2(n548), .Z(n549) );
  and2 U712 ( .A1(n601), .A2(n630), .Z(n571) );
  inv1 U713 ( .I(r), .ZN(n930) );
  inv1 U716 ( .I(n846), .ZN(n844) );
  or2 U717 ( .A1(n512), .A2(n887), .Z(n890) );
  inv1 U724 ( .I(n894), .ZN(n892) );
  or2 U735 ( .A1(n938), .A2(n937), .Z(n939) );
  inv1f U736 ( .I(n1012), .ZN(n540) );
  inv1 U740 ( .I(n1004), .ZN(n536) );
  inv1 U741 ( .I(n942), .ZN(n1023) );
  inv1 U742 ( .I(n966), .ZN(n1027) );
  or2 U743 ( .A1(n719), .A2(n718), .Z(n966) );
  or2 U744 ( .A1(n820), .A2(n819), .Z(n970) );
  inv1f U745 ( .I(t), .ZN(n937) );
  inv1f U748 ( .I(n511), .ZN(n917) );
  or2f U749 ( .A1(n960), .A2(n1000), .Z(n947) );
  or2f U757 ( .A1(n681), .A2(n680), .Z(n684) );
  or2f U758 ( .A1(n785), .A2(n784), .Z(n788) );
  or2f U762 ( .A1(n814), .A2(n813), .Z(n817) );
  inv1 U763 ( .I(n970), .ZN(n1025) );
  inv1 U764 ( .I(n1025), .ZN(n1026) );
  inv1 U769 ( .I(n1023), .ZN(n1024) );
  and2f U770 ( .A1(n933), .A2(t), .Z(n693) );
  inv1f U772 ( .I(h), .ZN(n516) );
  or2f U773 ( .A1(n1013), .A2(n537), .Z(n1006) );
  or2f U774 ( .A1(n936), .A2(n541), .Z(n938) );
  inv1f U778 ( .I(n540), .ZN(n541) );
  and2f U779 ( .A1(s), .A2(n937), .Z(n692) );
  inv1 U795 ( .I(n1027), .ZN(n1028) );
  or2f U798 ( .A1(n995), .A2(n968), .Z(n972) );
  inv1f U808 ( .I(n607), .ZN(n604) );
  or2f U809 ( .A1(n960), .A2(n541), .Z(n963) );
  or2f U810 ( .A1(n960), .A2(n537), .Z(n952) );
  or2f U832 ( .A1(n960), .A2(n533), .Z(n957) );
  or2f U835 ( .A1(n578), .A2(n577), .Z(n1000) );
  and2f U836 ( .A1(n917), .A2(n1000), .Z(n918) );
  or2 U868 ( .A1(n541), .A2(n1000), .Z(n850) );
  or2f U870 ( .A1(n988), .A2(n537), .Z(n980) );
  or2f U872 ( .A1(n988), .A2(n533), .Z(n985) );
  and2f U873 ( .A1(n821), .A2(n997), .Z(n824) );
  or2f U884 ( .A1(n695), .A2(n694), .Z(n698) );
  and2f U891 ( .A1(n930), .A2(q), .Z(n694) );
  or2f U893 ( .A1(n969), .A2(n966), .Z(n924) );
  or2f U895 ( .A1(n609), .A2(n608), .Z(n612) );
  or2f U897 ( .A1(n520), .A2(n533), .Z(n934) );
  and2f U898 ( .A1(n822), .A2(n924), .Z(n823) );
  or2f U899 ( .A1(n729), .A2(n728), .Z(n802) );
  and2f U900 ( .A1(n818), .A2(n817), .Z(n819) );
  or2f U901 ( .A1(n529), .A2(n533), .Z(n1010) );
  and2f U902 ( .A1(n597), .A2(n596), .Z(n598) );
  inv1f U903 ( .I(n595), .ZN(n597) );
  or2f U904 ( .A1(n843), .A2(n1024), .Z(n846) );
  or2f U905 ( .A1(n843), .A2(n1028), .Z(n830) );
  or2f U906 ( .A1(n891), .A2(n1024), .Z(n894) );
  or2f U907 ( .A1(n891), .A2(n1028), .Z(n879) );
  and2f U908 ( .A1(n642), .A2(n641), .Z(n646) );
  inv1 U913 ( .I(n643), .ZN(n641) );
  or2f U916 ( .A1(n633), .A2(n632), .Z(n636) );
  and2f U918 ( .A1(n630), .A2(n528), .Z(n633) );
  or2f U921 ( .A1(n936), .A2(n1000), .Z(n928) );
  or2f U923 ( .A1(n926), .A2(n925), .Z(n936) );
  or2f U924 ( .A1(n995), .A2(n941), .Z(n944) );
  or2f U928 ( .A1(n560), .A2(n559), .Z(n601) );
  and2f U930 ( .A1(n558), .A2(n557), .Z(n559) );
  and2f U931 ( .A1(n671), .A2(n670), .Z(n675) );
  or2f U932 ( .A1(n662), .A2(n661), .Z(n665) );
  and2f U933 ( .A1(n660), .A2(n528), .Z(n661) );
  or2f U937 ( .A1(n988), .A2(n541), .Z(n991) );
  and2f U938 ( .A1(r), .A2(n927), .Z(n695) );
  or2f U942 ( .A1(n867), .A2(n1024), .Z(n869) );
  or2f U943 ( .A1(n867), .A2(n1028), .Z(n854) );
  and2f U947 ( .A1(n966), .A2(n969), .Z(n821) );
  or2f U948 ( .A1(n912), .A2(n1024), .Z(n914) );
  or2f U955 ( .A1(n912), .A2(n1028), .Z(n901) );
  or2f U956 ( .A1(n520), .A2(n537), .Z(n931) );
  or2f U957 ( .A1(n926), .A2(n925), .Z(n520) );
  and2f U962 ( .A1(n595), .A2(n594), .Z(n599) );
  inv1f U965 ( .I(n596), .ZN(n594) );
  or2f U967 ( .A1(n995), .A2(n994), .Z(n999) );
  and2f U968 ( .A1(n613), .A2(n612), .Z(n614) );
  or2f U969 ( .A1(n843), .A2(n1026), .Z(n835) );
  or2f U972 ( .A1(n891), .A2(n1026), .Z(n884) );
  or2f U973 ( .A1(n867), .A2(n1026), .Z(n859) );
  or2f U978 ( .A1(n912), .A2(n1026), .Z(n905) );
  and2f U979 ( .A1(n970), .A2(n942), .Z(n822) );
  or2f U980 ( .A1(n646), .A2(n645), .Z(n1012) );
  and2f U984 ( .A1(n636), .A2(n635), .Z(n640) );
  or2f U985 ( .A1(n599), .A2(n598), .Z(n658) );
  or2f U989 ( .A1(n598), .A2(n599), .Z(n513) );
  or2f U990 ( .A1(n675), .A2(n674), .Z(n1004) );
  and2f U994 ( .A1(n665), .A2(n664), .Z(n669) );
  inv1f U995 ( .I(n665), .ZN(n667) );
  or2f U999 ( .A1(n867), .A2(n969), .Z(n864) );
  or2f U1001 ( .A1(n851), .A2(n898), .Z(n867) );
  or2f U1003 ( .A1(n755), .A2(n754), .Z(n969) );
  and2f U1004 ( .A1(n751), .A2(n750), .Z(n755) );
  or2f U1005 ( .A1(n640), .A2(n639), .Z(n643) );
  and2f U1006 ( .A1(n638), .A2(n637), .Z(n639) );
  or2f U1007 ( .A1(n529), .A2(n541), .Z(n1015) );
  or2f U1009 ( .A1(n999), .A2(n998), .Z(n529) );
  or2f U1010 ( .A1(n301), .A2(n302), .Z(n299) );
  and2f U1013 ( .A1(m), .A2(n1020), .Z(n302) );
  and2f U1016 ( .A1(n298), .A2(n627), .Z(n628) );
  or2f U1019 ( .A1(n303), .A2(n304), .Z(n298) );
  or2f U1020 ( .A1(n944), .A2(n943), .Z(n960) );
  or2f U1024 ( .A1(n988), .A2(n1000), .Z(n975) );
  or2f U1026 ( .A1(n972), .A2(n971), .Z(n988) );
  and2f U1027 ( .A1(n611), .A2(n610), .Z(n615) );
  or2f U1028 ( .A1(n629), .A2(n628), .Z(n659) );
  or2f U1032 ( .A1(n843), .A2(n969), .Z(n840) );
  or2f U1033 ( .A1(n827), .A2(n826), .Z(n843) );
  or2f U1037 ( .A1(n536), .A2(n873), .Z(n826) );
  and2f U1038 ( .A1(n816), .A2(n815), .Z(n820) );
  or2f U1042 ( .A1(n912), .A2(n969), .Z(n909) );
  or2f U1043 ( .A1(n899), .A2(n898), .Z(n912) );
  or2f U1047 ( .A1(n701), .A2(n700), .Z(n738) );
  and2f U1049 ( .A1(n699), .A2(n698), .Z(n700) );
  or2f U1051 ( .A1(n873), .A2(n532), .Z(n898) );
  and2f U1052 ( .A1(n919), .A2(n541), .Z(n920) );
  or2f U1053 ( .A1(n995), .A2(n1025), .Z(n926) );
  and2f U1057 ( .A1(n685), .A2(n684), .Z(n686) );
  inv1f U1058 ( .I(n825), .ZN(n873) );
  or2f U1062 ( .A1(n824), .A2(n823), .Z(n825) );
  or2f U1063 ( .A1(n876), .A2(n875), .Z(n891) );
  or2f U1067 ( .A1(n540), .A2(n873), .Z(n875) );
  and2f U1068 ( .A1(n536), .A2(n540), .Z(n511) );
  or2f U1072 ( .A1(n669), .A2(n668), .Z(n672) );
  and2f U1074 ( .A1(n667), .A2(n666), .Z(n668) );
  or2f U1075 ( .A1(n1013), .A2(n1000), .Z(n1002) );
  or2f U1078 ( .A1(n999), .A2(n998), .Z(n1013) );
  or2f U1081 ( .A1(n922), .A2(n921), .Z(n923) );
  or2f U1084 ( .A1(n564), .A2(n563), .Z(n508) );
  or2f U1087 ( .A1(n570), .A2(n569), .Z(n631) );
  and2f U1088 ( .A1(n566), .A2(n565), .Z(n570) );
  or2f U1089 ( .A1(n570), .A2(n509), .Z(n510) );
  inv1f U1090 ( .I(n923), .ZN(n995) );
endmodule

