
module unreg ( k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, 
        s, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, a1, z0, y0, x0, 
        w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0 );
  input k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, q,
         p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0;
  wire   n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184;

  inv1 U109 ( .I(t), .ZN(n92) );
  and2 U111 ( .A1(d), .A2(n87), .Z(n97) );
  inv1 U112 ( .I(w), .ZN(n102) );
  inv1 U114 ( .I(s), .ZN(n94) );
  and2 U116 ( .A1(n102), .A2(n182), .Z(n96) );
  inv1 U118 ( .I(v), .ZN(n129) );
  inv1 U119 ( .I(u), .ZN(n175) );
  and2 U120 ( .A1(n129), .A2(n175), .Z(n98) );
  or2 U121 ( .A1(n99), .A2(n98), .Z(l0) );
  inv1 U123 ( .I(x), .ZN(n107) );
  and2 U124 ( .A1(n107), .A2(n88), .Z(n100) );
  or2 U125 ( .A1(n101), .A2(n100), .Z(n104) );
  and2 U126 ( .A1(n102), .A2(n175), .Z(n103) );
  or2 U127 ( .A1(n104), .A2(n103), .Z(m0) );
  inv1 U129 ( .I(y), .ZN(n112) );
  and2 U130 ( .A1(n112), .A2(n183), .Z(n105) );
  or2 U131 ( .A1(n106), .A2(n105), .Z(n109) );
  and2 U132 ( .A1(n107), .A2(n175), .Z(n108) );
  or2 U133 ( .A1(n109), .A2(n108), .Z(n0) );
  or2 U136 ( .A1(n111), .A2(n110), .Z(n114) );
  and2 U137 ( .A1(n112), .A2(n175), .Z(n113) );
  or2 U138 ( .A1(n114), .A2(n113), .Z(o0) );
  inv1 U140 ( .I(a0), .ZN(n121) );
  and2 U141 ( .A1(n121), .A2(n183), .Z(n115) );
  or2 U142 ( .A1(n116), .A2(n115), .Z(n118) );
  inv1 U143 ( .I(z), .ZN(n149) );
  and2 U144 ( .A1(n149), .A2(n175), .Z(n117) );
  or2 U145 ( .A1(n118), .A2(n117), .Z(p0) );
  and2 U146 ( .A1(g), .A2(n87), .Z(n120) );
  inv1 U147 ( .I(b0), .ZN(n126) );
  and2 U150 ( .A1(n121), .A2(n175), .Z(n122) );
  or2 U151 ( .A1(n123), .A2(n122), .Z(q0) );
  inv1 U153 ( .I(c0), .ZN(n132) );
  or2 U155 ( .A1(n125), .A2(n124), .Z(n128) );
  and2 U156 ( .A1(n126), .A2(n175), .Z(n127) );
  or2 U157 ( .A1(n128), .A2(n127), .Z(r0) );
  and2 U159 ( .A1(n129), .A2(n88), .Z(n130) );
  or2 U160 ( .A1(n131), .A2(n130), .Z(n134) );
  and2 U161 ( .A1(n132), .A2(n175), .Z(n133) );
  or2 U162 ( .A1(n134), .A2(n133), .Z(s0) );
  inv1 U164 ( .I(e0), .ZN(n141) );
  or2 U166 ( .A1(n136), .A2(n135), .Z(n138) );
  inv1 U167 ( .I(d0), .ZN(n172) );
  and2 U168 ( .A1(n172), .A2(n175), .Z(n137) );
  or2 U169 ( .A1(n138), .A2(n137), .Z(t0) );
  inv1 U171 ( .I(f0), .ZN(n146) );
  and2 U172 ( .A1(n146), .A2(n88), .Z(n139) );
  or2 U173 ( .A1(n140), .A2(n139), .Z(n143) );
  and2 U174 ( .A1(n141), .A2(n175), .Z(n142) );
  or2 U175 ( .A1(n143), .A2(n142), .Z(u0) );
  inv1 U177 ( .I(g0), .ZN(n152) );
  and2 U178 ( .A1(n152), .A2(n182), .Z(n144) );
  or2 U179 ( .A1(n145), .A2(n144), .Z(n148) );
  and2 U180 ( .A1(n146), .A2(n175), .Z(n147) );
  or2 U181 ( .A1(n148), .A2(n147), .Z(v0) );
  and2 U183 ( .A1(n149), .A2(n183), .Z(n150) );
  or2 U184 ( .A1(n151), .A2(n150), .Z(n154) );
  and2 U185 ( .A1(n152), .A2(n175), .Z(n153) );
  or2 U186 ( .A1(n154), .A2(n153), .Z(w0) );
  and2 U187 ( .A1(p), .A2(n87), .Z(n156) );
  inv1 U188 ( .I(i0), .ZN(n162) );
  and2 U189 ( .A1(n162), .A2(n182), .Z(n155) );
  inv1 U191 ( .I(h0), .ZN(n157) );
  and2 U192 ( .A1(n157), .A2(n175), .Z(n158) );
  or2 U193 ( .A1(n159), .A2(n158), .Z(x0) );
  inv1 U195 ( .I(j0), .ZN(n167) );
  and2 U196 ( .A1(n167), .A2(n88), .Z(n160) );
  or2 U197 ( .A1(n161), .A2(n160), .Z(n164) );
  and2 U198 ( .A1(n162), .A2(n175), .Z(n163) );
  or2 U199 ( .A1(n164), .A2(n163), .Z(y0) );
  inv1 U201 ( .I(k0), .ZN(n176) );
  and2 U202 ( .A1(n176), .A2(n183), .Z(n165) );
  or2 U203 ( .A1(n166), .A2(n165), .Z(n169) );
  and2 U204 ( .A1(n167), .A2(n175), .Z(n168) );
  or2 U205 ( .A1(n169), .A2(n168), .Z(z0) );
  and2 U206 ( .A1(m), .A2(n87), .Z(n174) );
  and2 U207 ( .A1(n172), .A2(n182), .Z(n173) );
  and2 U209 ( .A1(n176), .A2(n175), .Z(n177) );
  or2 U210 ( .A1(n178), .A2(n177), .Z(a1) );
  inv1 U103 ( .I(s), .ZN(n91) );
  and2 U104 ( .A1(q), .A2(n171), .Z(n110) );
  and2 U105 ( .A1(n126), .A2(n171), .Z(n119) );
  and2 U106 ( .A1(n132), .A2(n171), .Z(n124) );
  and2 U107 ( .A1(n141), .A2(n171), .Z(n135) );
  and2f U108 ( .A1(u), .A2(t), .Z(n179) );
  and2f U110 ( .A1(l), .A2(n170), .Z(n136) );
  and2f U113 ( .A1(k), .A2(n170), .Z(n140) );
  and2f U115 ( .A1(h), .A2(n170), .Z(n116) );
  and2f U117 ( .A1(i), .A2(n90), .Z(n151) );
  and2f U122 ( .A1(e), .A2(n90), .Z(n131) );
  and2f U128 ( .A1(j), .A2(n90), .Z(n145) );
  and2f U134 ( .A1(o), .A2(n184), .Z(n161) );
  and2f U135 ( .A1(a), .A2(n184), .Z(n111) );
  and2f U139 ( .A1(f), .A2(n184), .Z(n125) );
  and2f U148 ( .A1(n), .A2(n89), .Z(n166) );
  and2f U149 ( .A1(b), .A2(n89), .Z(n106) );
  and2f U152 ( .A1(c), .A2(n89), .Z(n101) );
  or2f U154 ( .A1(n97), .A2(n96), .Z(n99) );
  or2f U158 ( .A1(n120), .A2(n119), .Z(n123) );
  or2f U163 ( .A1(n156), .A2(n155), .Z(n159) );
  or2f U165 ( .A1(n174), .A2(n173), .Z(n178) );
  and2f U170 ( .A1(u), .A2(n91), .Z(n181) );
  and2f U176 ( .A1(u), .A2(n91), .Z(n180) );
  and2f U182 ( .A1(n179), .A2(n94), .Z(n171) );
  and2f U190 ( .A1(n181), .A2(n92), .Z(n170) );
  and2f U194 ( .A1(n180), .A2(n92), .Z(n90) );
  and2f U200 ( .A1(n181), .A2(n92), .Z(n89) );
  and2f U208 ( .A1(n95), .A2(n94), .Z(n183) );
  and2f U211 ( .A1(n179), .A2(n94), .Z(n182) );
  and2f U212 ( .A1(u), .A2(t), .Z(n95) );
  and2f U213 ( .A1(n95), .A2(n94), .Z(n88) );
  and2f U214 ( .A1(n180), .A2(n92), .Z(n184) );
  and2f U215 ( .A1(u), .A2(n91), .Z(n93) );
  and2f U216 ( .A1(n93), .A2(n92), .Z(n87) );
endmodule

