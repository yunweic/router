
module vda ( q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, d1, c1, b1, a1, 
        z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, 
        h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r );
  input q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0,
         m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u,
         t, s, r;
  wire   n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n224, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519;

  or2f U1 ( .A1(n21), .A2(n22), .Z(y0) );
  or2f U2 ( .A1(n25), .A2(n496), .Z(n22) );
  or2f U10 ( .A1(n35), .A2(n36), .Z(v0) );
  or2f U13 ( .A1(n40), .A2(n41), .Z(n25) );
  or2f U14 ( .A1(n476), .A2(n43), .Z(n41) );
  or2f U19 ( .A1(n488), .A2(n52), .Z(n47) );
  or2f U20 ( .A1(n466), .A2(n53), .Z(n52) );
  or2f U23 ( .A1(n58), .A2(n59), .Z(n466) );
  or2f U24 ( .A1(n60), .A2(n61), .Z(n59) );
  or2f U25 ( .A1(n62), .A2(n63), .Z(t0) );
  or2f U26 ( .A1(n64), .A2(n37), .Z(n63) );
  or2f U33 ( .A1(n73), .A2(n74), .Z(r0) );
  or2f U34 ( .A1(n75), .A2(n76), .Z(n74) );
  or2f U35 ( .A1(n23), .A2(n499), .Z(n76) );
  or2f U38 ( .A1(n34), .A2(n79), .Z(n61) );
  or2f U40 ( .A1(n81), .A2(n82), .Z(r) );
  or2f U42 ( .A1(n488), .A2(n83), .Z(n81) );
  or2f U43 ( .A1(n85), .A2(n502), .Z(n83) );
  or2f U45 ( .A1(n86), .A2(n87), .Z(n85) );
  or2f U46 ( .A1(n42), .A2(n57), .Z(n87) );
  or2f U48 ( .A1(n89), .A2(n90), .Z(n88) );
  or2f U50 ( .A1(n463), .A2(n93), .Z(n92) );
  or2f U57 ( .A1(n54), .A2(n30), .Z(n458) );
  or2f U59 ( .A1(n49), .A2(n101), .Z(n43) );
  or2f U61 ( .A1(n104), .A2(n105), .Z(o0) );
  or2f U62 ( .A1(n64), .A2(n106), .Z(n105) );
  or2f U63 ( .A1(n107), .A2(n108), .Z(n64) );
  or2f U64 ( .A1(n109), .A2(n110), .Z(n108) );
  or2f U72 ( .A1(n118), .A2(n119), .Z(m0) );
  or2f U79 ( .A1(n23), .A2(n91), .Z(n32) );
  or2f U80 ( .A1(n124), .A2(n125), .Z(n23) );
  or2f U82 ( .A1(n117), .A2(n127), .Z(l0) );
  or2f U84 ( .A1(n128), .A2(n111), .Z(n90) );
  or2f U85 ( .A1(n474), .A2(n96), .Z(n117) );
  or2f U88 ( .A1(n86), .A2(n132), .Z(n96) );
  or2f U93 ( .A1(n135), .A2(n136), .Z(k0) );
  or2f U94 ( .A1(n482), .A2(n453), .Z(n136) );
  or2f U96 ( .A1(n515), .A2(n476), .Z(n138) );
  or2f U98 ( .A1(n141), .A2(n142), .Z(n140) );
  or2f U99 ( .A1(n26), .A2(n143), .Z(n142) );
  or2f U101 ( .A1(n146), .A2(n147), .Z(n139) );
  and2f U104 ( .A1(n467), .A2(n149), .Z(n124) );
  or2f U105 ( .A1(n150), .A2(n151), .Z(n42) );
  or2f U106 ( .A1(n152), .A2(n100), .Z(n151) );
  or2f U113 ( .A1(n158), .A2(n159), .Z(n157) );
  or2f U114 ( .A1(n160), .A2(n161), .Z(n159) );
  or2f U115 ( .A1(n38), .A2(n162), .Z(n161) );
  or2f U131 ( .A1(n183), .A2(n184), .Z(h0) );
  or2f U132 ( .A1(n185), .A2(n186), .Z(n184) );
  or2f U135 ( .A1(n189), .A2(n190), .Z(n160) );
  or2f U136 ( .A1(n191), .A2(n192), .Z(n190) );
  and2f U154 ( .A1(c), .A2(n215), .Z(n111) );
  and2f U155 ( .A1(n170), .A2(n216), .Z(n215) );
  or2f U159 ( .A1(n220), .A2(n221), .Z(g0) );
  and2f U175 ( .A1(n239), .A2(e), .Z(n93) );
  and2f U177 ( .A1(n242), .A2(n243), .Z(n241) );
  or2f U179 ( .A1(n246), .A2(n247), .Z(n245) );
  or2f U182 ( .A1(n251), .A2(n252), .Z(n250) );
  or2f U183 ( .A1(n253), .A2(n254), .Z(n252) );
  or2f U184 ( .A1(n49), .A2(n255), .Z(n251) );
  or2f U185 ( .A1(n256), .A2(n257), .Z(n49) );
  and2f U190 ( .A1(n262), .A2(n210), .Z(n261) );
  and2f U198 ( .A1(n262), .A2(i), .Z(n144) );
  or2f U226 ( .A1(n295), .A2(n296), .Z(e0) );
  or2f U227 ( .A1(n297), .A2(n298), .Z(n296) );
  or2f U228 ( .A1(n226), .A2(n299), .Z(n298) );
  or2f U236 ( .A1(n209), .A2(n309), .Z(n300) );
  or2f U237 ( .A1(n456), .A2(n310), .Z(n309) );
  or2f U241 ( .A1(n314), .A2(n315), .Z(n187) );
  or2f U242 ( .A1(n316), .A2(n317), .Z(n315) );
  and2f U248 ( .A1(n494), .A2(n325), .Z(n322) );
  and2f U251 ( .A1(n327), .A2(n328), .Z(n320) );
  and2f U254 ( .A1(n332), .A2(h), .Z(n327) );
  or2f U261 ( .A1(n227), .A2(n337), .Z(n143) );
  or2f U262 ( .A1(n44), .A2(n229), .Z(n337) );
  and2f U264 ( .A1(n232), .A2(n313), .Z(n304) );
  and2f U266 ( .A1(n313), .A2(n281), .Z(n338) );
  or2f U271 ( .A1(n342), .A2(n343), .Z(n314) );
  and2f U282 ( .A1(n170), .A2(n271), .Z(n262) );
  and2f U294 ( .A1(n170), .A2(n334), .Z(n267) );
  or2f U299 ( .A1(n361), .A2(n362), .Z(n360) );
  or2f U300 ( .A1(n224), .A2(n248), .Z(n362) );
  or2f U307 ( .A1(n366), .A2(n367), .Z(n224) );
  or2f U308 ( .A1(n368), .A2(n369), .Z(n367) );
  or2f U310 ( .A1(n370), .A2(n371), .Z(n71) );
  and2f U314 ( .A1(n180), .A2(n238), .Z(n375) );
  and2f U318 ( .A1(n334), .A2(n378), .Z(n370) );
  or2f U319 ( .A1(n379), .A2(n380), .Z(n378) );
  and2f U321 ( .A1(n381), .A2(n382), .Z(n379) );
  or2f U322 ( .A1(n383), .A2(n305), .Z(n381) );
  and2f U323 ( .A1(n384), .A2(m), .Z(n383) );
  and2f U324 ( .A1(n230), .A2(n210), .Z(n384) );
  and2f U329 ( .A1(n171), .A2(n356), .Z(n216) );
  or2f U342 ( .A1(n72), .A2(n394), .Z(n391) );
  or2f U343 ( .A1(n145), .A2(n100), .Z(n394) );
  or2f U351 ( .A1(n253), .A2(n401), .Z(n361) );
  or2f U352 ( .A1(n402), .A2(n162), .Z(n401) );
  or2f U353 ( .A1(n403), .A2(n404), .Z(n162) );
  or2f U364 ( .A1(n409), .A2(n410), .Z(n408) );
  or2f U367 ( .A1(n411), .A2(n412), .Z(n409) );
  and2f U370 ( .A1(n395), .A2(c), .Z(n413) );
  or2f U374 ( .A1(n285), .A2(n44), .Z(n415) );
  inv1f U375 ( .I(n416), .ZN(n285) );
  or2f U376 ( .A1(n330), .A2(n417), .Z(n416) );
  or2f U377 ( .A1(n411), .A2(n382), .Z(n417) );
  inv1f U379 ( .I(n377), .ZN(n411) );
  and2f U380 ( .A1(n468), .A2(n418), .Z(n377) );
  and2f U381 ( .A1(n210), .A2(n334), .Z(n418) );
  or2f U383 ( .A1(n168), .A2(n242), .Z(n330) );
  or2f U384 ( .A1(b), .A2(n336), .Z(n242) );
  and2f U387 ( .A1(n334), .A2(n364), .Z(n44) );
  and2f U406 ( .A1(n238), .A2(n428), .Z(n152) );
  and2f U410 ( .A1(n169), .A2(q), .Z(n356) );
  and2f U413 ( .A1(l), .A2(o), .Z(n238) );
  and2f U416 ( .A1(n171), .A2(n232), .Z(n180) );
  and2f U421 ( .A1(h), .A2(n430), .Z(n310) );
  and2f U422 ( .A1(n334), .A2(n305), .Z(n430) );
  and2f U423 ( .A1(n431), .A2(n), .Z(n334) );
  and2f U425 ( .A1(n400), .A2(l), .Z(n270) );
  or2f U427 ( .A1(n39), .A2(n461), .Z(n50) );
  and2f U431 ( .A1(n169), .A2(n433), .Z(n396) );
  and2f U432 ( .A1(n434), .A2(g), .Z(n39) );
  or2f U433 ( .A1(n435), .A2(n436), .Z(n434) );
  and2f U435 ( .A1(n230), .A2(n282), .Z(n305) );
  and2f U436 ( .A1(n467), .A2(m), .Z(n282) );
  inv1f U439 ( .I(n), .ZN(n169) );
  and2f U441 ( .A1(n), .A2(n433), .Z(n271) );
  and2f U443 ( .A1(n294), .A2(p), .Z(n202) );
  and2f U446 ( .A1(n174), .A2(n170), .Z(n281) );
  and2f U447 ( .A1(n308), .A2(n400), .Z(n170) );
  inv1f U448 ( .I(o), .ZN(n400) );
  and2f U451 ( .A1(n294), .A2(n148), .Z(n171) );
  inv1f U453 ( .I(m), .ZN(n294) );
  buf0 U454 ( .I(n465), .Z(t) );
  buf0 U455 ( .I(n466), .Z(u) );
  buf0 U456 ( .I(n465), .Z(w) );
  buf0 U457 ( .I(n465), .Z(x) );
  buf0 U458 ( .I(n464), .Z(y) );
  buf0 U459 ( .I(n463), .Z(z) );
  buf0 U460 ( .I(n462), .Z(a0) );
  buf0 U461 ( .I(n461), .Z(b0) );
  buf0 U462 ( .I(n460), .Z(c0) );
  buf0 U463 ( .I(n459), .Z(j0) );
  buf0 U464 ( .I(n458), .Z(p0) );
  buf0 U465 ( .I(n457), .Z(z0) );
  buf0 U466 ( .I(n456), .Z(a1) );
  buf0 U467 ( .I(n455), .Z(b1) );
  buf0 U468 ( .I(n454), .Z(c1) );
  buf0 U469 ( .I(n453), .Z(d1) );
  or2f U470 ( .A1(n488), .A2(n39), .Z(n137) );
  inv1f U471 ( .I(p), .ZN(n148) );
  inv1f U472 ( .I(q), .ZN(n431) );
  and2f U473 ( .A1(q), .A2(n), .Z(n174) );
  or2f U474 ( .A1(n179), .A2(n344), .Z(n343) );
  or2f U475 ( .A1(n60), .A2(n34), .Z(n346) );
  and2f U476 ( .A1(n294), .A2(n230), .Z(n365) );
  or2f U477 ( .A1(n133), .A2(n89), .Z(n201) );
  and2f U478 ( .A1(n232), .A2(n238), .Z(n292) );
  and2f U479 ( .A1(n396), .A2(n238), .Z(n425) );
  and2f U480 ( .A1(n232), .A2(n170), .Z(n203) );
  and2f U481 ( .A1(n243), .A2(n395), .Z(n100) );
  and2f U482 ( .A1(n170), .A2(n396), .Z(n243) );
  or2 U483 ( .A1(n144), .A2(n145), .Z(n26) );
  and2 U484 ( .A1(n322), .A2(n323), .Z(n321) );
  and2 U485 ( .A1(n230), .A2(n271), .Z(n435) );
  inv1 U486 ( .I(n495), .ZN(n468) );
  or2 U487 ( .A1(n501), .A2(n45), .Z(n268) );
  or2 U488 ( .A1(n150), .A2(n204), .Z(n199) );
  or2 U489 ( .A1(n241), .A2(n240), .Z(n239) );
  or2 U490 ( .A1(n420), .A2(n421), .Z(n253) );
  and2 U491 ( .A1(k), .A2(n426), .Z(n344) );
  or2 U492 ( .A1(n391), .A2(n392), .Z(n366) );
  and2 U493 ( .A1(g), .A2(n425), .Z(n51) );
  and2 U494 ( .A1(n261), .A2(d), .Z(n256) );
  or2 U495 ( .A1(n92), .A2(n490), .Z(n502) );
  or2 U496 ( .A1(n91), .A2(n92), .Z(n84) );
  or2 U497 ( .A1(n460), .A2(n461), .Z(n512) );
  and2 U498 ( .A1(a), .A2(n292), .Z(n291) );
  or2 U499 ( .A1(n106), .A2(n160), .Z(n188) );
  and2 U500 ( .A1(n262), .A2(n348), .Z(n53) );
  inv1 U501 ( .I(n214), .ZN(n510) );
  or2 U502 ( .A1(n475), .A2(n515), .Z(n54) );
  and2 U503 ( .A1(n236), .A2(n203), .Z(n60) );
  or2 U504 ( .A1(n112), .A2(n113), .Z(n107) );
  or2 U505 ( .A1(n124), .A2(n485), .Z(n496) );
  or2 U506 ( .A1(n156), .A2(n157), .Z(i0) );
  or2 U507 ( .A1(n30), .A2(n31), .Z(x0) );
  inv1 U508 ( .I(p), .ZN(n467) );
  or2 U509 ( .A1(n80), .A2(n56), .Z(n79) );
  and2f U510 ( .A1(n173), .A2(n174), .Z(n80) );
  and2f U511 ( .A1(n294), .A2(n472), .Z(n433) );
  and2f U512 ( .A1(n468), .A2(n418), .Z(n469) );
  or2f U513 ( .A1(n), .A2(q), .Z(n470) );
  inv1f U514 ( .I(n470), .ZN(n232) );
  and2f U515 ( .A1(n171), .A2(n232), .Z(n471) );
  or2f U516 ( .A1(n460), .A2(n102), .Z(n58) );
  or2 U517 ( .A1(n511), .A2(n512), .Z(n462) );
  and2 U518 ( .A1(n434), .A2(g), .Z(n511) );
  and2 U519 ( .A1(n329), .A2(n), .Z(n328) );
  and2 U520 ( .A1(n330), .A2(n331), .Z(n329) );
  inv1 U521 ( .I(m), .ZN(n484) );
  or2 U522 ( .A1(n60), .A2(n53), .Z(n172) );
  and2 U523 ( .A1(n243), .A2(b), .Z(n287) );
  or2 U524 ( .A1(n462), .A2(n46), .Z(n132) );
  or2 U525 ( .A1(n34), .A2(n43), .Z(n99) );
  inv1 U526 ( .I(l), .ZN(n308) );
  and2 U527 ( .A1(g), .A2(n325), .Z(n258) );
  and2 U528 ( .A1(a), .A2(n375), .Z(n240) );
  or2 U529 ( .A1(n372), .A2(n373), .Z(n371) );
  and2 U530 ( .A1(n376), .A2(n469), .Z(n372) );
  and2 U531 ( .A1(n375), .A2(n480), .Z(n373) );
  or2 U532 ( .A1(n300), .A2(n301), .Z(n254) );
  or2 U533 ( .A1(n263), .A2(n264), .Z(n249) );
  and2 U534 ( .A1(n322), .A2(n323), .Z(n492) );
  or2 U535 ( .A1(n320), .A2(n321), .Z(n319) );
  or2 U536 ( .A1(n199), .A2(n200), .Z(n189) );
  or2 U537 ( .A1(n272), .A2(n415), .Z(n403) );
  or2 U538 ( .A1(n152), .A2(n58), .Z(n277) );
  or2 U539 ( .A1(n413), .A2(n288), .Z(n412) );
  and2 U540 ( .A1(n270), .A2(n356), .Z(n397) );
  and2 U541 ( .A1(n270), .A2(n282), .Z(n364) );
  and2 U542 ( .A1(n396), .A2(n432), .Z(n461) );
  or2 U543 ( .A1(n115), .A2(n66), .Z(n141) );
  or2 U544 ( .A1(n80), .A2(n172), .Z(n103) );
  and2 U545 ( .A1(n267), .A2(n335), .Z(n78) );
  or2 U546 ( .A1(n91), .A2(n38), .Z(n499) );
  or2 U547 ( .A1(n67), .A2(n88), .Z(n57) );
  or2 U548 ( .A1(n359), .A2(n360), .Z(d0) );
  or2 U549 ( .A1(n244), .A2(n245), .Z(f0) );
  or2 U550 ( .A1(n98), .A2(n99), .Z(n94) );
  or2 U551 ( .A1(n458), .A2(n67), .Z(s0) );
  and2 U552 ( .A1(p), .A2(q), .Z(n472) );
  buf0 U553 ( .I(n49), .Z(n473) );
  or2 U554 ( .A1(n56), .A2(n43), .Z(n30) );
  and2 U555 ( .A1(n326), .A2(n304), .Z(n229) );
  and2 U556 ( .A1(n326), .A2(e), .Z(n332) );
  or2f U557 ( .A1(n67), .A2(n405), .Z(n404) );
  or2f U558 ( .A1(n198), .A2(n268), .Z(n263) );
  or2 U559 ( .A1(n516), .A2(n50), .Z(n110) );
  or2 U560 ( .A1(n193), .A2(n194), .Z(n192) );
  and2f U561 ( .A1(n243), .A2(n487), .Z(n193) );
  or2 U562 ( .A1(n497), .A2(n27), .Z(n474) );
  or2 U563 ( .A1(n85), .A2(n84), .Z(n465) );
  or2 U564 ( .A1(n96), .A2(n486), .Z(n130) );
  or2 U565 ( .A1(n94), .A2(n95), .Z(q0) );
  or2 U566 ( .A1(n126), .A2(n89), .Z(n421) );
  or2f U567 ( .A1(n126), .A2(n149), .Z(n204) );
  or2 U568 ( .A1(n476), .A2(n137), .Z(n475) );
  or2 U569 ( .A1(n482), .A2(n55), .Z(u0) );
  or2f U570 ( .A1(n150), .A2(n151), .Z(n476) );
  or2f U571 ( .A1(n241), .A2(n479), .Z(n477) );
  and2f U572 ( .A1(n477), .A2(n478), .Z(n125) );
  or2 U573 ( .A1(n126), .A2(e), .Z(n478) );
  or2 U574 ( .A1(n240), .A2(n126), .Z(n479) );
  and2 U575 ( .A1(a), .A2(n374), .Z(n480) );
  and2 U576 ( .A1(n232), .A2(n305), .Z(n436) );
  or2 U577 ( .A1(n23), .A2(n481), .Z(w0) );
  and2f U578 ( .A1(n238), .A2(n271), .Z(n56) );
  or2f U579 ( .A1(n197), .A2(n198), .Z(n196) );
  or2 U580 ( .A1(n91), .A2(n33), .Z(n481) );
  or2f U581 ( .A1(n138), .A2(n137), .Z(n482) );
  or2f U582 ( .A1(n148), .A2(n484), .Z(n483) );
  inv1 U583 ( .I(n483), .ZN(n236) );
  and2 U584 ( .A1(n236), .A2(n397), .Z(n145) );
  and2 U585 ( .A1(n236), .A2(n338), .Z(n227) );
  and2 U586 ( .A1(n232), .A2(n326), .Z(n325) );
  and2 U587 ( .A1(n326), .A2(n333), .Z(n177) );
  or2 U588 ( .A1(n125), .A2(n516), .Z(n485) );
  or2 U589 ( .A1(n27), .A2(n106), .Z(n486) );
  and2 U590 ( .A1(b), .A2(n286), .Z(n487) );
  and2 U591 ( .A1(g), .A2(n425), .Z(n488) );
  and2f U592 ( .A1(n356), .A2(n238), .Z(n385) );
  or2f U593 ( .A1(n32), .A2(n122), .Z(n118) );
  or2f U594 ( .A1(n370), .A2(n489), .Z(n369) );
  or2f U595 ( .A1(n371), .A2(n37), .Z(n489) );
  or2 U596 ( .A1(n91), .A2(n39), .Z(n490) );
  and2 U597 ( .A1(n286), .A2(n287), .Z(n491) );
  or2f U598 ( .A1(n492), .A2(n493), .Z(n255) );
  or2 U599 ( .A1(n318), .A2(n320), .Z(n493) );
  and2 U600 ( .A1(g), .A2(n168), .Z(n494) );
  or2f U601 ( .A1(n503), .A2(n483), .Z(n495) );
  inv1f U602 ( .I(n495), .ZN(n326) );
  and2 U603 ( .A1(n258), .A2(n259), .Z(n257) );
  or2f U604 ( .A1(n227), .A2(n228), .Z(n38) );
  or2f U605 ( .A1(n463), .A2(n229), .Z(n228) );
  or2f U606 ( .A1(n140), .A2(n139), .Z(n86) );
  or2f U607 ( .A1(n140), .A2(n139), .Z(n515) );
  or2 U608 ( .A1(n106), .A2(n129), .Z(n497) );
  or2 U609 ( .A1(n130), .A2(n498), .Z(n0) );
  or2 U610 ( .A1(n129), .A2(n116), .Z(n498) );
  and2f U611 ( .A1(n239), .A2(e), .Z(n500) );
  and2f U612 ( .A1(n230), .A2(n396), .Z(n426) );
  and2f U613 ( .A1(n313), .A2(n396), .Z(n428) );
  and2f U614 ( .A1(n270), .A2(n396), .Z(n456) );
  or2f U615 ( .A1(n187), .A2(n188), .Z(n186) );
  or2f U616 ( .A1(n317), .A2(n316), .Z(n517) );
  or2f U617 ( .A1(n319), .A2(n519), .Z(n317) );
  or2f U618 ( .A1(n32), .A2(n516), .Z(n31) );
  or2 U619 ( .A1(n500), .A2(n114), .Z(n112) );
  and2f U620 ( .A1(n262), .A2(i), .Z(n501) );
  or2 U621 ( .A1(n96), .A2(n97), .Z(n95) );
  or2f U622 ( .A1(l), .A2(n504), .Z(n503) );
  inv1f U623 ( .I(n503), .ZN(n230) );
  inv1f U624 ( .I(o), .ZN(n504) );
  or2 U625 ( .A1(n250), .A2(n249), .Z(n505) );
  or2f U626 ( .A1(n505), .A2(n506), .Z(n221) );
  or2f U627 ( .A1(n224), .A2(n222), .Z(n506) );
  or2f U628 ( .A1(n251), .A2(n252), .Z(n507) );
  or2f U629 ( .A1(n507), .A2(n508), .Z(n247) );
  or2 U630 ( .A1(n248), .A2(n249), .Z(n508) );
  and2f U631 ( .A1(n408), .A2(n510), .Z(n509) );
  inv1f U632 ( .I(n509), .ZN(n67) );
  inv1 U633 ( .I(n408), .ZN(n114) );
  or2f U634 ( .A1(n39), .A2(n25), .Z(n35) );
  or2f U635 ( .A1(n53), .A2(n60), .Z(n513) );
  or2f U636 ( .A1(n513), .A2(n514), .Z(n101) );
  or2 U637 ( .A1(n102), .A2(n80), .Z(n514) );
  or2 U638 ( .A1(n501), .A2(n145), .Z(n516) );
  and2f U639 ( .A1(n202), .A2(n292), .Z(n89) );
  or2f U640 ( .A1(n517), .A2(n518), .Z(n299) );
  or2 U641 ( .A1(n254), .A2(n314), .Z(n518) );
  or2 U642 ( .A1(n318), .A2(n143), .Z(n519) );
  and2 U643 ( .A1(n236), .A2(n390), .Z(n351) );
  and2 U644 ( .A1(l), .A2(n232), .Z(n390) );
  inv1 U645 ( .I(e), .ZN(n288) );
  or2 U646 ( .A1(n347), .A2(n53), .Z(n226) );
  and2 U647 ( .A1(n350), .A2(n174), .Z(n347) );
  and2 U648 ( .A1(n171), .A2(l), .Z(n350) );
  or2 U649 ( .A1(n45), .A2(n123), .Z(n147) );
  and2 U650 ( .A1(n270), .A2(n471), .Z(n420) );
  and2 U651 ( .A1(n171), .A2(n267), .Z(n46) );
  or2 U652 ( .A1(c), .A2(n260), .Z(n259) );
  and2 U653 ( .A1(n210), .A2(n324), .Z(n323) );
  and2 U654 ( .A1(g), .A2(n236), .Z(n306) );
  and2 U655 ( .A1(n174), .A2(n308), .Z(n307) );
  and2 U656 ( .A1(n304), .A2(n305), .Z(n303) );
  inv1 U657 ( .I(j), .ZN(n331) );
  inv1 U658 ( .I(h), .ZN(n382) );
  inv1 U659 ( .I(k), .ZN(n324) );
  or2 U660 ( .A1(n206), .A2(n363), .Z(n248) );
  or2 U661 ( .A1(n149), .A2(n453), .Z(n363) );
  and2 U662 ( .A1(n173), .A2(n334), .Z(n272) );
  and2 U663 ( .A1(n288), .A2(f), .Z(n286) );
  and2 U664 ( .A1(n270), .A2(n202), .Z(n341) );
  or2 U665 ( .A1(n265), .A2(n266), .Z(n264) );
  or2 U666 ( .A1(n155), .A2(n197), .Z(n392) );
  or2 U667 ( .A1(n453), .A2(n346), .Z(n342) );
  and2 U668 ( .A1(n334), .A2(n345), .Z(n179) );
  and2 U669 ( .A1(n171), .A2(o), .Z(n345) );
  and2 U670 ( .A1(n202), .A2(n203), .Z(n128) );
  and2 U671 ( .A1(f), .A2(n414), .Z(n395) );
  inv1 U672 ( .I(b), .ZN(n414) );
  and2 U673 ( .A1(n230), .A2(n231), .Z(n219) );
  and2 U674 ( .A1(n202), .A2(n232), .Z(n231) );
  or2 U675 ( .A1(n51), .A2(n461), .Z(n275) );
  and2 U676 ( .A1(n232), .A2(n341), .Z(n214) );
  and2 U677 ( .A1(n238), .A2(n216), .Z(n123) );
  and2 U678 ( .A1(n230), .A2(n216), .Z(n91) );
  and2 U679 ( .A1(n267), .A2(n279), .Z(n133) );
  and2 U680 ( .A1(n202), .A2(f), .Z(n279) );
  and2 U681 ( .A1(n471), .A2(n170), .Z(n70) );
  and2 U682 ( .A1(n398), .A2(n399), .Z(n72) );
  and2 U683 ( .A1(n400), .A2(n336), .Z(n398) );
  and2 U684 ( .A1(n288), .A2(n396), .Z(n399) );
  or2 U685 ( .A1(n457), .A2(n152), .Z(n427) );
  and2 U686 ( .A1(n419), .A2(n236), .Z(n402) );
  and2 U687 ( .A1(n334), .A2(n400), .Z(n419) );
  or2 U688 ( .A1(n344), .A2(n424), .Z(n423) );
  or2 U689 ( .A1(n488), .A2(n456), .Z(n424) );
  and2 U690 ( .A1(n282), .A2(n267), .Z(n164) );
  or2 U691 ( .A1(n351), .A2(n352), .Z(n297) );
  or2 U692 ( .A1(n285), .A2(n353), .Z(n352) );
  or2 U693 ( .A1(n357), .A2(n358), .Z(n354) );
  or2 U694 ( .A1(n152), .A2(n56), .Z(n358) );
  or2 U695 ( .A1(n39), .A2(n145), .Z(n357) );
  and2 U696 ( .A1(n290), .A2(n291), .Z(n195) );
  and2 U697 ( .A1(f), .A2(n293), .Z(n290) );
  and2 U698 ( .A1(n294), .A2(n288), .Z(n293) );
  or2 U699 ( .A1(n179), .A2(n164), .Z(n289) );
  or2 U700 ( .A1(n272), .A2(n75), .Z(n246) );
  or2 U701 ( .A1(n491), .A2(n285), .Z(n284) );
  and2 U702 ( .A1(n334), .A2(n341), .Z(n235) );
  and2 U703 ( .A1(n236), .A2(n237), .Z(n194) );
  and2 U704 ( .A1(n169), .A2(n238), .Z(n237) );
  or2 U705 ( .A1(n38), .A2(n226), .Z(n222) );
  or2 U706 ( .A1(n93), .A2(n91), .Z(n233) );
  or2 U707 ( .A1(n123), .A2(n214), .Z(n213) );
  or2 U708 ( .A1(n473), .A2(n205), .Z(n185) );
  or2 U709 ( .A1(n206), .A2(n207), .Z(n205) );
  and2 U710 ( .A1(n208), .A2(n209), .Z(n207) );
  and2 U711 ( .A1(n168), .A2(n210), .Z(n208) );
  or2 U712 ( .A1(n217), .A2(n218), .Z(n211) );
  or2 U713 ( .A1(n460), .A2(n91), .Z(n218) );
  or2 U714 ( .A1(n454), .A2(n219), .Z(n217) );
  and2 U715 ( .A1(n334), .A2(i), .Z(n333) );
  or2 U716 ( .A1(n70), .A2(n179), .Z(n178) );
  or2 U717 ( .A1(n103), .A2(n163), .Z(n158) );
  or2 U718 ( .A1(n164), .A2(n165), .Z(n163) );
  and2 U719 ( .A1(n166), .A2(n167), .Z(n165) );
  and2 U720 ( .A1(n168), .A2(n169), .Z(n167) );
  or2 U721 ( .A1(n181), .A2(n182), .Z(n175) );
  or2 U722 ( .A1(n66), .A2(n46), .Z(n182) );
  or2 U723 ( .A1(n45), .A2(n100), .Z(n181) );
  or2 U724 ( .A1(n123), .A2(n66), .Z(n122) );
  or2 U725 ( .A1(n476), .A2(n121), .Z(n116) );
  or2 U726 ( .A1(n454), .A2(n488), .Z(n121) );
  or2 U727 ( .A1(n453), .A2(n134), .Z(n129) );
  or2 U728 ( .A1(n89), .A2(n456), .Z(n134) );
  and2 U729 ( .A1(n356), .A2(n326), .Z(n115) );
  or2 U730 ( .A1(n457), .A2(n455), .Z(n106) );
  or2 U731 ( .A1(n71), .A2(n154), .Z(n459) );
  or2 U732 ( .A1(n70), .A2(n155), .Z(n154) );
  or2 U733 ( .A1(n219), .A2(n29), .Z(n463) );
  or2 U734 ( .A1(n27), .A2(n67), .Z(n97) );
  and2 U735 ( .A1(n210), .A2(n349), .Z(n348) );
  inv1 U736 ( .I(d), .ZN(n349) );
  and2 U737 ( .A1(n336), .A2(n202), .Z(n335) );
  or2 U738 ( .A1(n273), .A2(n274), .Z(n75) );
  or2 U739 ( .A1(n277), .A2(n278), .Z(n273) );
  or2 U740 ( .A1(n275), .A2(n276), .Z(n274) );
  or2 U741 ( .A1(n150), .A2(n133), .Z(n278) );
  and2 U742 ( .A1(n282), .A2(n203), .Z(n66) );
  or2 U743 ( .A1(n111), .A2(n46), .Z(n109) );
  or2 U744 ( .A1(n44), .A2(n45), .Z(n40) );
  or2 U745 ( .A1(n123), .A2(n34), .Z(n37) );
  and2 U746 ( .A1(n282), .A2(n385), .Z(n34) );
  and2 U747 ( .A1(n230), .A2(n471), .Z(n29) );
  and2 U748 ( .A1(n171), .A2(n281), .Z(n460) );
  or2 U749 ( .A1(n133), .A2(n78), .Z(n27) );
  and2 U750 ( .A1(n173), .A2(n356), .Z(n457) );
  and2 U751 ( .A1(j), .A2(n310), .Z(n455) );
  or2 U752 ( .A1(n429), .A2(n420), .Z(n454) );
  and2 U753 ( .A1(n326), .A2(n174), .Z(n429) );
  and2 U754 ( .A1(n174), .A2(n364), .Z(n453) );
  inv1 U755 ( .I(a), .ZN(n389) );
  or2 U756 ( .A1(n78), .A2(n177), .Z(n318) );
  and2 U757 ( .A1(n270), .A2(n271), .Z(n198) );
  and2 U758 ( .A1(n236), .A2(n406), .Z(n265) );
  and2 U759 ( .A1(n356), .A2(n170), .Z(n406) );
  and2 U760 ( .A1(n267), .A2(n236), .Z(n266) );
  and2 U761 ( .A1(n356), .A2(n364), .Z(n197) );
  or2 U762 ( .A1(n351), .A2(n386), .Z(n368) );
  and2 U763 ( .A1(n387), .A2(n388), .Z(n386) );
  and2 U764 ( .A1(n169), .A2(n467), .Z(n388) );
  and2 U765 ( .A1(n238), .A2(n389), .Z(n387) );
  or2 U766 ( .A1(n235), .A2(n339), .Z(n316) );
  and2 U767 ( .A1(n340), .A2(n282), .Z(n339) );
  and2 U768 ( .A1(n170), .A2(q), .Z(n340) );
  or2 U769 ( .A1(n195), .A2(n196), .Z(n191) );
  or2 U770 ( .A1(n128), .A2(n201), .Z(n200) );
  or2 U771 ( .A1(n353), .A2(n265), .Z(n405) );
  or2 U772 ( .A1(n126), .A2(n124), .Z(n146) );
  inv1 U773 ( .I(g), .ZN(n313) );
  and2 U774 ( .A1(n281), .A2(n282), .Z(n102) );
  and2 U775 ( .A1(n334), .A2(n365), .Z(n149) );
  and2 U776 ( .A1(n330), .A2(n288), .Z(n376) );
  and2 U777 ( .A1(n238), .A2(n202), .Z(n380) );
  and2 U778 ( .A1(n288), .A2(n336), .Z(n374) );
  or2 U779 ( .A1(n302), .A2(n303), .Z(n301) );
  and2 U780 ( .A1(n306), .A2(n307), .Z(n302) );
  and2 U781 ( .A1(m), .A2(n407), .Z(n353) );
  and2 U782 ( .A1(n270), .A2(n232), .Z(n407) );
  and2 U783 ( .A1(n311), .A2(n312), .Z(n209) );
  and2 U784 ( .A1(n313), .A2(p), .Z(n311) );
  and2 U785 ( .A1(n230), .A2(n174), .Z(n312) );
  and2 U786 ( .A1(n356), .A2(n305), .Z(n206) );
  inv1 U787 ( .I(c), .ZN(n168) );
  and2 U788 ( .A1(n170), .A2(n171), .Z(n166) );
  and2 U789 ( .A1(n334), .A2(n393), .Z(n155) );
  and2 U790 ( .A1(n238), .A2(n282), .Z(n393) );
  inv1 U791 ( .I(i), .ZN(n210) );
  inv1 U792 ( .I(f), .ZN(n336) );
  and2 U793 ( .A1(n174), .A2(n280), .Z(n150) );
  and2 U794 ( .A1(n171), .A2(n230), .Z(n280) );
  or2 U795 ( .A1(n115), .A2(n46), .Z(n276) );
  or2 U796 ( .A1(n382), .A2(n331), .Z(n410) );
  or2 U797 ( .A1(n29), .A2(n89), .Z(n113) );
  or2 U798 ( .A1(k), .A2(i), .Z(n260) );
  and2 U799 ( .A1(n236), .A2(n269), .Z(n45) );
  and2 U800 ( .A1(n270), .A2(n174), .Z(n269) );
  and2 U801 ( .A1(n292), .A2(n282), .Z(n126) );
  and2 U802 ( .A1(n270), .A2(n171), .Z(n173) );
  or2 U803 ( .A1(n47), .A2(n48), .Z(n464) );
  or2 U804 ( .A1(n49), .A2(n50), .Z(n48) );
  and2 U805 ( .A1(n324), .A2(n230), .Z(n432) );
  or2 U806 ( .A1(n46), .A2(n27), .Z(n82) );
  or2 U807 ( .A1(n456), .A2(n72), .Z(n68) );
  or2 U808 ( .A1(n70), .A2(n71), .Z(n69) );
  or2 U809 ( .A1(n464), .A2(n46), .Z(v) );
  or2 U810 ( .A1(n422), .A2(n423), .Z(n359) );
  or2 U811 ( .A1(n56), .A2(n427), .Z(n422) );
  or2 U812 ( .A1(n354), .A2(n355), .Z(n295) );
  or2 U813 ( .A1(n164), .A2(n141), .Z(n355) );
  or2 U814 ( .A1(n283), .A2(n284), .Z(n244) );
  or2 U815 ( .A1(n195), .A2(n289), .Z(n283) );
  or2 U816 ( .A1(n233), .A2(n234), .Z(n220) );
  or2 U817 ( .A1(n194), .A2(n235), .Z(n234) );
  or2 U818 ( .A1(n211), .A2(n212), .Z(n183) );
  or2 U819 ( .A1(n111), .A2(n213), .Z(n212) );
  or2 U820 ( .A1(n175), .A2(n176), .Z(n156) );
  or2 U821 ( .A1(n177), .A2(n178), .Z(n176) );
  or2 U822 ( .A1(n455), .A2(n153), .Z(n135) );
  or2 U823 ( .A1(n459), .A2(n454), .Z(n153) );
  or2 U824 ( .A1(n463), .A2(n90), .Z(n127) );
  or2 U825 ( .A1(n116), .A2(n120), .Z(n119) );
  or2 U826 ( .A1(n90), .A2(n38), .Z(n120) );
  or2 U827 ( .A1(n459), .A2(n115), .Z(n104) );
  or2 U828 ( .A1(n463), .A2(n100), .Z(n98) );
  or2 U829 ( .A1(n61), .A2(n77), .Z(n73) );
  or2 U830 ( .A1(n53), .A2(n78), .Z(n77) );
  or2 U831 ( .A1(n473), .A2(n65), .Z(n62) );
  or2 U832 ( .A1(n60), .A2(n66), .Z(n65) );
  or2 U833 ( .A1(n56), .A2(n57), .Z(n55) );
  or2 U834 ( .A1(n37), .A2(n38), .Z(n36) );
  or2 U835 ( .A1(n34), .A2(n516), .Z(n33) );
  or2 U836 ( .A1(n27), .A2(n28), .Z(n21) );
  or2 U837 ( .A1(n29), .A2(n460), .Z(n28) );
  or2 U838 ( .A1(n68), .A2(n69), .Z(s) );
endmodule

