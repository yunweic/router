
module alu4_cl ( j, i, h, g, f, e, d, c, b, a, p, o, n, m, l, k );
  input j, i, h, g, f, e, d, c, b, a;
  output p, o, n, m, l, k;
  wire   n741, n60, n61, n62, n93, n124, n126, n147, n148, n291, n292, n295,
         n300, n301, n302, n303, n315, n316, n328, n330, n335, n346, n347,
         n348, n352, n402, n403, n407, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n456, n458, n459, n460, n461, n462, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n503, n504, n505, n506, n507, n508, n512, n513, n514,
         n515, n517, n518, n519, n521, n522, n523, n526, n527, n528, n529,
         n530, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n574, n576, n579, n580, n581,
         n582, n584, n585, n586, n587, n588, n589, n590, n591, n595, n597,
         n598, n599, n602, n603, n604, n605, n606, n607, n608, n610, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n632, n633, n634, n635,
         n636, n637, n638, n639, n642, n643, n644, n645, n646, n647, n648,
         n649, n654, n655, n656, n659, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n701,
         n702, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n735, n736, n738,
         n739, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837;

  or2f U9 ( .A1(n61), .A2(n62), .Z(n60) );
  or2f U214 ( .A1(n291), .A2(n292), .Z(k) );
  and2f U255 ( .A1(n330), .A2(j), .Z(n291) );
  and2f U274 ( .A1(n346), .A2(n347), .Z(n335) );
  or2f U280 ( .A1(n352), .A2(h), .Z(n346) );
  or2f U364 ( .A1(n795), .A2(h), .Z(n403) );
  buf0 U366 ( .I(n741), .Z(m) );
  buf0 U367 ( .I(n739), .Z(n) );
  or2 U370 ( .A1(n830), .A2(n806), .Z(n470) );
  or2 U371 ( .A1(n830), .A2(g), .Z(n645) );
  or2 U375 ( .A1(n793), .A2(h), .Z(n705) );
  or2 U376 ( .A1(n770), .A2(n821), .Z(n570) );
  or2 U377 ( .A1(n402), .A2(n643), .Z(n458) );
  and2 U378 ( .A1(n643), .A2(n619), .Z(n467) );
  or2 U379 ( .A1(n758), .A2(n619), .Z(n620) );
  or2 U380 ( .A1(n619), .A2(g), .Z(n460) );
  or2 U381 ( .A1(n832), .A2(a), .Z(n454) );
  and2f U390 ( .A1(n699), .A2(n819), .Z(n732) );
  and2 U392 ( .A1(n626), .A2(n708), .Z(n627) );
  or2 U394 ( .A1(n708), .A2(b), .Z(n713) );
  and2 U395 ( .A1(n743), .A2(n701), .Z(n702) );
  and2 U396 ( .A1(n663), .A2(n743), .Z(n544) );
  and2 U397 ( .A1(n490), .A2(n556), .Z(n487) );
  and2 U398 ( .A1(b), .A2(n744), .Z(n561) );
  and2 U399 ( .A1(b), .A2(n708), .Z(n709) );
  or2 U400 ( .A1(n708), .A2(n664), .Z(n665) );
  and2 U401 ( .A1(n807), .A2(n708), .Z(n603) );
  or2 U402 ( .A1(n708), .A2(n643), .Z(n644) );
  or2 U403 ( .A1(n830), .A2(n663), .Z(n604) );
  or2 U406 ( .A1(n744), .A2(n643), .Z(n581) );
  or2 U408 ( .A1(n708), .A2(n752), .Z(n547) );
  inv1f U417 ( .I(f), .ZN(n668) );
  inv1f U419 ( .I(g), .ZN(n663) );
  inv1f U421 ( .I(n415), .ZN(n673) );
  and2f U422 ( .A1(n802), .A2(n673), .Z(n418) );
  and2f U425 ( .A1(n490), .A2(n416), .Z(n417) );
  or2f U426 ( .A1(n418), .A2(n417), .Z(n422) );
  and2f U430 ( .A1(h), .A2(n808), .Z(n419) );
  and2f U431 ( .A1(n663), .A2(n419), .Z(n420) );
  or2f U433 ( .A1(n420), .A2(n690), .Z(n421) );
  or2f U434 ( .A1(n422), .A2(n421), .Z(n423) );
  and2f U435 ( .A1(n424), .A2(n423), .Z(n432) );
  or2f U437 ( .A1(f), .A2(n563), .Z(n569) );
  or2f U440 ( .A1(n425), .A2(j), .Z(n428) );
  and2f U441 ( .A1(n403), .A2(n773), .Z(n426) );
  or2f U442 ( .A1(n426), .A2(n690), .Z(n427) );
  and2f U443 ( .A1(n427), .A2(n428), .Z(n430) );
  inv1f U445 ( .I(n643), .ZN(n714) );
  and2f U446 ( .A1(n556), .A2(n714), .Z(n429) );
  or2f U447 ( .A1(n430), .A2(n429), .Z(n533) );
  or2f U449 ( .A1(n432), .A2(n431), .Z(n441) );
  and2f U453 ( .A1(n633), .A2(n433), .Z(n439) );
  or2f U456 ( .A1(n436), .A2(n821), .Z(n437) );
  and2f U459 ( .A1(n534), .A2(n480), .Z(n438) );
  or2f U460 ( .A1(n439), .A2(n438), .Z(n440) );
  or2f U461 ( .A1(n441), .A2(n440), .Z(n642) );
  or2f U472 ( .A1(n796), .A2(n446), .Z(n447) );
  or2f U473 ( .A1(n781), .A2(n447), .Z(n448) );
  and2f U474 ( .A1(n556), .A2(n448), .Z(n449) );
  and2f U475 ( .A1(n820), .A2(n829), .Z(n451) );
  or2f U476 ( .A1(n452), .A2(n451), .Z(n465) );
  or2f U494 ( .A1(n466), .A2(n832), .Z(n469) );
  and2f U496 ( .A1(n469), .A2(n468), .Z(n472) );
  and2f U499 ( .A1(n472), .A2(n471), .Z(n473) );
  and2f U501 ( .A1(n783), .A2(n346), .Z(n475) );
  or2f U502 ( .A1(n792), .A2(n690), .Z(n477) );
  or2f U543 ( .A1(n824), .A2(g), .Z(n508) );
  inv1f U544 ( .I(n508), .ZN(n571) );
  and2f U555 ( .A1(n556), .A2(n662), .Z(n515) );
  or2f U557 ( .A1(n515), .A2(n799), .Z(n517) );
  and2f U558 ( .A1(n518), .A2(n517), .Z(n519) );
  or2f U566 ( .A1(n802), .A2(n668), .Z(n526) );
  and2f U567 ( .A1(n527), .A2(n526), .Z(n528) );
  or2f U568 ( .A1(n528), .A2(n529), .Z(n530) );
  and2f U571 ( .A1(n533), .A2(n682), .Z(n539) );
  and2f U572 ( .A1(n534), .A2(n720), .Z(n537) );
  and2f U573 ( .A1(h), .A2(n571), .Z(n535) );
  or2f U575 ( .A1(n537), .A2(n536), .Z(n538) );
  or2f U576 ( .A1(n539), .A2(n538), .Z(n540) );
  or2f U577 ( .A1(n541), .A2(n540), .Z(n708) );
  or2f U587 ( .A1(n625), .A2(n549), .Z(n550) );
  or2f U590 ( .A1(n708), .A2(n551), .Z(n552) );
  or2f U592 ( .A1(n678), .A2(n553), .Z(n554) );
  or2f U593 ( .A1(n554), .A2(n683), .Z(n555) );
  and2f U594 ( .A1(n555), .A2(n556), .Z(n559) );
  or2f U596 ( .A1(n559), .A2(n558), .Z(n698) );
  and2f U608 ( .A1(n610), .A2(n681), .Z(n572) );
  and2f U620 ( .A1(n402), .A2(n585), .Z(n588) );
  and2f U622 ( .A1(n597), .A2(n586), .Z(n587) );
  or2f U623 ( .A1(n588), .A2(n587), .Z(n589) );
  and2f U631 ( .A1(b), .A2(n602), .Z(n607) );
  or2f U634 ( .A1(n607), .A2(n606), .Z(n608) );
  and2f U638 ( .A1(n613), .A2(n695), .Z(n614) );
  or2f U639 ( .A1(n614), .A2(g), .Z(n615) );
  or2f U640 ( .A1(n616), .A2(n615), .Z(n624) );
  or2f U666 ( .A1(n655), .A2(n656), .Z(n699) );
  or2f U696 ( .A1(n702), .A2(n60), .Z(n707) );
  inv1 U362 ( .I(n748), .ZN(n742) );
  and2f U363 ( .A1(n762), .A2(n763), .Z(n602) );
  or2 U365 ( .A1(n754), .A2(e), .Z(n752) );
  inv1f U368 ( .I(g), .ZN(n795) );
  inv1 U369 ( .I(n772), .ZN(n579) );
  inv1 U372 ( .I(n751), .ZN(n434) );
  inv1 U373 ( .I(e), .ZN(n563) );
  or2 U374 ( .A1(n522), .A2(j), .Z(n523) );
  inv1 U382 ( .I(a), .ZN(n803) );
  inv1 U383 ( .I(b), .ZN(n626) );
  inv1 U384 ( .I(n809), .ZN(n613) );
  inv1 U385 ( .I(n624), .ZN(n774) );
  or2 U386 ( .A1(n828), .A2(n654), .Z(n769) );
  inv1f U387 ( .I(n465), .ZN(n749) );
  and2f U388 ( .A1(n714), .A2(n698), .Z(n585) );
  inv1f U389 ( .I(e), .ZN(n822) );
  or2f U391 ( .A1(n441), .A2(n440), .Z(n766) );
  inv1f U393 ( .I(n610), .ZN(n744) );
  inv1f U404 ( .I(n698), .ZN(n610) );
  inv1f U405 ( .I(n708), .ZN(n625) );
  inv1 U407 ( .I(n582), .ZN(n704) );
  or2 U409 ( .A1(n581), .A2(n402), .Z(n582) );
  inv1 U410 ( .I(n523), .ZN(n529) );
  or2 U411 ( .A1(n414), .A2(j), .Z(n424) );
  and2 U412 ( .A1(n557), .A2(n713), .Z(n558) );
  or2 U413 ( .A1(n705), .A2(n704), .Z(n706) );
  or2 U414 ( .A1(g), .A2(b), .Z(n522) );
  inv1 U415 ( .I(n794), .ZN(n425) );
  inv1 U416 ( .I(n413), .ZN(n414) );
  or2 U418 ( .A1(n412), .A2(n411), .Z(n413) );
  or2 U420 ( .A1(g), .A2(e), .Z(n412) );
  or2 U423 ( .A1(h), .A2(a), .Z(n411) );
  inv1 U424 ( .I(n437), .ZN(n534) );
  and2 U427 ( .A1(n435), .A2(n434), .Z(n436) );
  or2 U428 ( .A1(h), .A2(j), .Z(n435) );
  inv1 U429 ( .I(c), .ZN(n490) );
  and2 U432 ( .A1(g), .A2(a), .Z(n797) );
  inv1 U436 ( .I(n798), .ZN(n453) );
  inv1 U438 ( .I(n403), .ZN(n556) );
  and2 U439 ( .A1(n714), .A2(n535), .Z(n536) );
  or2 U444 ( .A1(n694), .A2(n512), .Z(n518) );
  inv1 U448 ( .I(n513), .ZN(n664) );
  inv1 U450 ( .I(n514), .ZN(n662) );
  or2 U451 ( .A1(b), .A2(n682), .Z(n514) );
  or2 U452 ( .A1(n473), .A2(n721), .Z(n474) );
  inv1 U454 ( .I(n550), .ZN(n683) );
  inv1 U455 ( .I(d), .ZN(n826) );
  inv1 U457 ( .I(b), .ZN(n825) );
  or2 U458 ( .A1(n561), .A2(n765), .Z(n562) );
  inv1 U462 ( .I(n623), .ZN(n810) );
  inv1 U463 ( .I(n639), .ZN(n811) );
  inv1 U464 ( .I(n612), .ZN(n616) );
  and2 U465 ( .A1(n574), .A2(n820), .Z(n580) );
  and2 U466 ( .A1(g), .A2(n812), .Z(n787) );
  or2 U467 ( .A1(n590), .A2(n589), .Z(n591) );
  or2 U468 ( .A1(b), .A2(d), .Z(n720) );
  inv1 U469 ( .I(n780), .ZN(n782) );
  or2 U470 ( .A1(n832), .A2(n749), .Z(n695) );
  or2 U471 ( .A1(a), .A2(c), .Z(n480) );
  inv1 U477 ( .I(n720), .ZN(n694) );
  inv1 U478 ( .I(i), .ZN(n746) );
  or2 U479 ( .A1(n730), .A2(n729), .Z(n731) );
  and2 U480 ( .A1(n728), .A2(n727), .Z(n730) );
  or2 U481 ( .A1(n707), .A2(n706), .Z(n728) );
  and2 U482 ( .A1(n659), .A2(n819), .Z(n756) );
  inv1 U483 ( .I(n625), .ZN(n743) );
  or2 U484 ( .A1(n475), .A2(n818), .Z(n800) );
  and2 U485 ( .A1(n766), .A2(n782), .Z(n781) );
  inv1 U486 ( .I(n552), .ZN(n678) );
  inv1 U487 ( .I(a), .ZN(n806) );
  or2 U488 ( .A1(n805), .A2(n806), .Z(n804) );
  or2 U489 ( .A1(f), .A2(e), .Z(n551) );
  inv1 U490 ( .I(n551), .ZN(n633) );
  inv1 U491 ( .I(n800), .ZN(n819) );
  or2f U492 ( .A1(n746), .A2(n747), .Z(n745) );
  inv1f U493 ( .I(n477), .ZN(n747) );
  or2f U495 ( .A1(n749), .A2(n619), .Z(n748) );
  or2f U497 ( .A1(n836), .A2(n758), .Z(n576) );
  or2 U498 ( .A1(n775), .A2(n654), .Z(n750) );
  inv1 U500 ( .I(d), .ZN(n682) );
  and2 U503 ( .A1(g), .A2(j), .Z(n751) );
  inv1 U504 ( .I(j), .ZN(n690) );
  inv1 U505 ( .I(n820), .ZN(n821) );
  or2f U506 ( .A1(n754), .A2(e), .Z(n753) );
  inv1f U507 ( .I(n753), .ZN(n773) );
  inv1f U508 ( .I(f), .ZN(n754) );
  or2 U509 ( .A1(n793), .A2(n576), .Z(n574) );
  and2 U510 ( .A1(n576), .A2(n793), .Z(n772) );
  buf0 U511 ( .I(n817), .Z(n755) );
  inv1 U512 ( .I(n837), .ZN(n659) );
  or2f U513 ( .A1(n757), .A2(n756), .Z(l) );
  or2f U514 ( .A1(n661), .A2(n693), .Z(n757) );
  buf0 U515 ( .I(n625), .Z(n758) );
  and2f U516 ( .A1(n837), .A2(n800), .Z(n661) );
  and2 U517 ( .A1(n597), .A2(n610), .Z(n598) );
  and2f U518 ( .A1(n761), .A2(n767), .Z(n759) );
  or2f U519 ( .A1(n759), .A2(n760), .Z(n837) );
  and2 U520 ( .A1(j), .A2(n656), .Z(n760) );
  and2f U521 ( .A1(n768), .A2(j), .Z(n761) );
  or2f U522 ( .A1(n598), .A2(n764), .Z(n762) );
  or2 U523 ( .A1(n663), .A2(n633), .Z(n763) );
  or2f U524 ( .A1(n599), .A2(n663), .Z(n764) );
  and2f U525 ( .A1(n831), .A2(a), .Z(n765) );
  inv1 U526 ( .I(n765), .ZN(n597) );
  or2f U527 ( .A1(n827), .A2(n769), .Z(n767) );
  and2f U528 ( .A1(n767), .A2(n768), .Z(n655) );
  or2f U529 ( .A1(n774), .A2(n750), .Z(n768) );
  inv1 U530 ( .I(n556), .ZN(n770) );
  or2f U531 ( .A1(n572), .A2(n571), .Z(n771) );
  inv1f U532 ( .I(n771), .ZN(n836) );
  and2f U533 ( .A1(n773), .A2(a), .Z(n416) );
  and2f U534 ( .A1(n490), .A2(n533), .Z(n431) );
  inv1 U535 ( .I(n832), .ZN(n402) );
  inv1 U536 ( .I(n831), .ZN(n832) );
  or2f U537 ( .A1(n649), .A2(n801), .Z(n775) );
  and2f U538 ( .A1(n830), .A2(n557), .Z(n450) );
  and2f U539 ( .A1(n459), .A2(n776), .Z(n352) );
  and2 U540 ( .A1(n458), .A2(n462), .Z(n776) );
  or2f U541 ( .A1(n732), .A2(n779), .Z(n777) );
  and2f U542 ( .A1(n777), .A2(n778), .Z(o) );
  or2 U545 ( .A1(n735), .A2(j), .Z(n778) );
  or2 U546 ( .A1(n731), .A2(n735), .Z(n779) );
  or2 U547 ( .A1(n806), .A2(n643), .Z(n780) );
  and2f U548 ( .A1(n474), .A2(n347), .Z(n783) );
  and2f U549 ( .A1(n832), .A2(n820), .Z(n784) );
  or2f U550 ( .A1(n784), .A2(n785), .Z(n798) );
  or2 U551 ( .A1(n766), .A2(n452), .Z(n785) );
  or2f U552 ( .A1(n753), .A2(n403), .Z(n415) );
  and2f U553 ( .A1(n788), .A2(n580), .Z(n786) );
  or2f U554 ( .A1(n786), .A2(n787), .Z(n827) );
  and2f U556 ( .A1(n579), .A2(g), .Z(n788) );
  inv1f U559 ( .I(n831), .ZN(n829) );
  or2f U560 ( .A1(n742), .A2(n791), .Z(n789) );
  and2f U561 ( .A1(n789), .A2(n790), .Z(n459) );
  or2 U562 ( .A1(n456), .A2(n454), .Z(n790) );
  or2f U563 ( .A1(n453), .A2(n456), .Z(n791) );
  and2f U564 ( .A1(n335), .A2(n474), .Z(n792) );
  inv1f U565 ( .I(n748), .ZN(n793) );
  or2f U569 ( .A1(n663), .A2(n569), .Z(n794) );
  and2f U570 ( .A1(n633), .A2(n805), .Z(n796) );
  inv1 U574 ( .I(n797), .ZN(n617) );
  or2f U578 ( .A1(n664), .A2(n802), .Z(n799) );
  or2f U579 ( .A1(n608), .A2(n595), .Z(n828) );
  or2 U580 ( .A1(n810), .A2(n811), .Z(n801) );
  and2f U581 ( .A1(n803), .A2(c), .Z(n802) );
  inv1 U582 ( .I(n802), .ZN(n512) );
  inv1 U583 ( .I(n804), .ZN(n407) );
  inv1f U584 ( .I(n642), .ZN(n805) );
  buf0 U585 ( .I(n773), .Z(n807) );
  and2f U586 ( .A1(a), .A2(c), .Z(n808) );
  inv1 U588 ( .I(n808), .ZN(n566) );
  and2f U589 ( .A1(n836), .A2(n744), .Z(n809) );
  inv1 U591 ( .I(n836), .ZN(n701) );
  or2 U595 ( .A1(n465), .A2(g), .Z(n466) );
  or2 U597 ( .A1(n613), .A2(n695), .Z(n612) );
  and2f U598 ( .A1(n745), .A2(n800), .Z(n330) );
  or2 U599 ( .A1(n704), .A2(n591), .Z(n812) );
  or2f U600 ( .A1(n403), .A2(n817), .Z(n813) );
  inv1f U601 ( .I(n813), .ZN(n527) );
  inv1 U602 ( .I(n755), .ZN(n739) );
  or2f U603 ( .A1(n571), .A2(n816), .Z(n814) );
  and2f U604 ( .A1(n814), .A2(n815), .Z(n521) );
  or2 U605 ( .A1(f), .A2(h), .Z(n815) );
  or2f U606 ( .A1(n797), .A2(f), .Z(n816) );
  or2f U607 ( .A1(n825), .A2(n826), .Z(n817) );
  or2 U609 ( .A1(n690), .A2(i), .Z(n818) );
  inv1 U610 ( .I(n569), .ZN(n820) );
  or2f U611 ( .A1(n668), .A2(n822), .Z(n643) );
  and2f U612 ( .A1(n765), .A2(n698), .Z(n599) );
  and2 U613 ( .A1(n822), .A2(n562), .Z(n62) );
  or2f U614 ( .A1(n530), .A2(n521), .Z(n834) );
  and2f U615 ( .A1(n823), .A2(n833), .Z(n541) );
  and2f U616 ( .A1(n834), .A2(n822), .Z(n823) );
  or2f U617 ( .A1(n825), .A2(n826), .Z(n824) );
  or2 U618 ( .A1(n626), .A2(d), .Z(n513) );
  buf0 U619 ( .I(n766), .Z(n830) );
  or2f U621 ( .A1(n450), .A2(n449), .Z(n831) );
  or2f U624 ( .A1(n530), .A2(n668), .Z(n835) );
  or2f U625 ( .A1(n519), .A2(n835), .Z(n833) );
  and2 U626 ( .A1(n808), .A2(n556), .Z(n433) );
  and2 U627 ( .A1(n619), .A2(n584), .Z(n590) );
  or2 U628 ( .A1(n729), .A2(n721), .Z(n647) );
  inv1 U629 ( .I(n565), .ZN(n719) );
  or2 U630 ( .A1(n564), .A2(n566), .Z(n565) );
  or2 U632 ( .A1(n628), .A2(n627), .Z(n629) );
  and2 U633 ( .A1(b), .A2(n625), .Z(n628) );
  or2 U635 ( .A1(n622), .A2(n643), .Z(n623) );
  and2 U636 ( .A1(n621), .A2(n620), .Z(n622) );
  and2 U637 ( .A1(n93), .A2(n618), .Z(n621) );
  or2 U641 ( .A1(n636), .A2(n635), .Z(n637) );
  inv1 U642 ( .I(n711), .ZN(n635) );
  and2 U643 ( .A1(n804), .A2(n630), .Z(n636) );
  inv1 U644 ( .I(n629), .ZN(n630) );
  and2 U645 ( .A1(n407), .A2(n629), .Z(n638) );
  inv1 U646 ( .I(n830), .ZN(n619) );
  or2 U647 ( .A1(f), .A2(n663), .Z(n456) );
  inv1 U648 ( .I(n501), .ZN(n461) );
  or2 U649 ( .A1(n714), .A2(n663), .Z(n632) );
  inv1 U650 ( .I(n547), .ZN(n584) );
  or2 U651 ( .A1(n634), .A2(n633), .Z(n711) );
  inv1 U652 ( .I(n632), .ZN(n634) );
  or2 U653 ( .A1(n821), .A2(g), .Z(n564) );
  inv1 U654 ( .I(n604), .ZN(n548) );
  inv1 U655 ( .I(n564), .ZN(n718) );
  and2 U656 ( .A1(n566), .A2(n718), .Z(n568) );
  or2 U657 ( .A1(n664), .A2(n662), .Z(n567) );
  or2 U658 ( .A1(n648), .A2(n647), .Z(n649) );
  or2 U659 ( .A1(n684), .A2(n683), .Z(n685) );
  and2 U660 ( .A1(n682), .A2(n681), .Z(n684) );
  or2 U661 ( .A1(n505), .A2(n504), .Z(n506) );
  or2 U662 ( .A1(n503), .A2(n781), .Z(n504) );
  or2 U663 ( .A1(n300), .A2(n295), .Z(n505) );
  and2 U664 ( .A1(n633), .A2(n501), .Z(n503) );
  inv1 U665 ( .I(n500), .ZN(n691) );
  or2 U667 ( .A1(n499), .A2(n328), .Z(n500) );
  or2 U668 ( .A1(h), .A2(g), .Z(n328) );
  or2 U669 ( .A1(n643), .A2(n690), .Z(n499) );
  inv1 U670 ( .I(n695), .ZN(n696) );
  inv1 U671 ( .I(n480), .ZN(n736) );
  or2 U672 ( .A1(n694), .A2(n739), .Z(n741) );
  and2 U673 ( .A1(n626), .A2(n633), .Z(n586) );
  or2 U674 ( .A1(n617), .A2(n626), .Z(n618) );
  and2 U675 ( .A1(n820), .A2(n808), .Z(n446) );
  and2 U676 ( .A1(n619), .A2(n718), .Z(n484) );
  and2 U677 ( .A1(n668), .A2(n667), .Z(n669) );
  or2 U678 ( .A1(n666), .A2(n665), .Z(n667) );
  and2 U679 ( .A1(n663), .A2(n662), .Z(n666) );
  and2 U680 ( .A1(d), .A2(n807), .Z(n670) );
  and2 U681 ( .A1(n663), .A2(n808), .Z(n452) );
  or2 U682 ( .A1(b), .A2(a), .Z(n93) );
  and2 U683 ( .A1(n694), .A2(n719), .Z(n648) );
  and2 U684 ( .A1(d), .A2(n718), .Z(n595) );
  or2 U685 ( .A1(n605), .A2(h), .Z(n606) );
  and2 U686 ( .A1(n604), .A2(n603), .Z(n605) );
  or2 U687 ( .A1(n638), .A2(n637), .Z(n639) );
  inv1 U688 ( .I(n460), .ZN(n479) );
  or2 U689 ( .A1(n486), .A2(n485), .Z(n489) );
  and2 U690 ( .A1(n807), .A2(n483), .Z(n486) );
  and2 U691 ( .A1(n721), .A2(n484), .Z(n485) );
  and2 U692 ( .A1(g), .A2(n808), .Z(n483) );
  and2 U693 ( .A1(n668), .A2(n487), .Z(n488) );
  and2 U694 ( .A1(n479), .A2(n478), .Z(n482) );
  and2 U695 ( .A1(c), .A2(n822), .Z(n478) );
  or2 U697 ( .A1(n496), .A2(n830), .Z(n498) );
  and2 U698 ( .A1(f), .A2(n808), .Z(n496) );
  and2 U699 ( .A1(c), .A2(n807), .Z(n497) );
  or2 U700 ( .A1(n493), .A2(n492), .Z(n495) );
  and2 U701 ( .A1(n668), .A2(n491), .Z(n492) );
  and2 U702 ( .A1(n802), .A2(n718), .Z(n493) );
  and2 U703 ( .A1(n490), .A2(a), .Z(n491) );
  or2 U704 ( .A1(n797), .A2(n633), .Z(n494) );
  or2 U705 ( .A1(n461), .A2(n752), .Z(n462) );
  or2 U706 ( .A1(g), .A2(n348), .Z(n347) );
  and2 U707 ( .A1(n470), .A2(n464), .Z(n348) );
  or2 U708 ( .A1(n512), .A2(n822), .Z(n464) );
  or2 U709 ( .A1(n632), .A2(n470), .Z(n471) );
  or2 U710 ( .A1(n467), .A2(a), .Z(n468) );
  or2 U711 ( .A1(n542), .A2(n633), .Z(n543) );
  and2 U712 ( .A1(d), .A2(n822), .Z(n542) );
  and2 U713 ( .A1(h), .A2(n672), .Z(n675) );
  or2 U714 ( .A1(n671), .A2(n124), .Z(n672) );
  and2 U715 ( .A1(g), .A2(b), .Z(n124) );
  or2 U716 ( .A1(n670), .A2(n669), .Z(n671) );
  and2 U717 ( .A1(n673), .A2(n694), .Z(n674) );
  and2 U718 ( .A1(n721), .A2(n545), .Z(n148) );
  and2 U719 ( .A1(n718), .A2(n758), .Z(n545) );
  and2 U720 ( .A1(n548), .A2(n584), .Z(n61) );
  and2 U721 ( .A1(n713), .A2(n712), .Z(n717) );
  and2 U722 ( .A1(n711), .A2(n710), .Z(n712) );
  or2 U723 ( .A1(n709), .A2(n407), .Z(n710) );
  and2 U724 ( .A1(n715), .A2(n714), .Z(n716) );
  inv1 U725 ( .I(n93), .ZN(n715) );
  or2 U726 ( .A1(n722), .A2(n721), .Z(n723) );
  and2 U727 ( .A1(n720), .A2(n719), .Z(n722) );
  inv1 U728 ( .I(h), .ZN(n721) );
  or2 U729 ( .A1(n479), .A2(n548), .Z(n501) );
  or2 U730 ( .A1(n315), .A2(n316), .Z(n295) );
  or2 U731 ( .A1(n482), .A2(n481), .Z(n315) );
  or2 U732 ( .A1(n489), .A2(n488), .Z(n316) );
  and2 U733 ( .A1(n736), .A2(n673), .Z(n481) );
  and2 U734 ( .A1(h), .A2(n301), .Z(n300) );
  or2 U735 ( .A1(n302), .A2(n303), .Z(n301) );
  or2 U736 ( .A1(n495), .A2(n494), .Z(n302) );
  or2 U737 ( .A1(n498), .A2(n497), .Z(n303) );
  and2 U738 ( .A1(g), .A2(n680), .Z(n686) );
  or2 U739 ( .A1(n679), .A2(n678), .Z(n680) );
  and2 U740 ( .A1(n807), .A2(n739), .Z(n679) );
  or2 U741 ( .A1(n676), .A2(n126), .Z(n688) );
  or2 U742 ( .A1(n147), .A2(n148), .Z(n126) );
  or2 U743 ( .A1(n675), .A2(n674), .Z(n676) );
  and2 U744 ( .A1(n544), .A2(n543), .Z(n147) );
  inv1 U745 ( .I(n570), .ZN(n681) );
  inv1 U746 ( .I(n646), .ZN(n729) );
  or2 U747 ( .A1(n645), .A2(n644), .Z(n646) );
  or2 U748 ( .A1(n726), .A2(n725), .Z(n727) );
  or2 U749 ( .A1(n724), .A2(n723), .Z(n725) );
  or2 U750 ( .A1(n717), .A2(n716), .Z(n726) );
  and2 U751 ( .A1(n718), .A2(n739), .Z(n724) );
  and2 U752 ( .A1(n739), .A2(n719), .Z(n656) );
  and2 U753 ( .A1(n568), .A2(n567), .Z(n654) );
  inv1 U754 ( .I(n443), .ZN(n557) );
  or2 U755 ( .A1(n442), .A2(n752), .Z(n443) );
  or2 U756 ( .A1(n721), .A2(n690), .Z(n442) );
  and2 U757 ( .A1(n820), .A2(n739), .Z(n553) );
  or2 U758 ( .A1(n643), .A2(n626), .Z(n549) );
  or2 U759 ( .A1(n692), .A2(n691), .Z(n693) );
  and2 U760 ( .A1(n690), .A2(n689), .Z(n692) );
  or2 U761 ( .A1(n688), .A2(n687), .Z(n689) );
  or2 U762 ( .A1(n686), .A2(n685), .Z(n687) );
  or2 U763 ( .A1(n691), .A2(n507), .Z(n292) );
  and2 U764 ( .A1(n690), .A2(n506), .Z(n507) );
  and2 U765 ( .A1(n744), .A2(n697), .Z(n735) );
  or2 U766 ( .A1(n696), .A2(n701), .Z(n697) );
  or2 U767 ( .A1(n808), .A2(n736), .Z(n738) );
  and2 U768 ( .A1(n741), .A2(n738), .Z(p) );
endmodule

