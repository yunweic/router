
module x3 ( h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, 
        q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, 
        y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, 
        g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, 
        o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, 
        w0, v0, u0, t0, s0, r0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, 
        c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, 
        f, e, d, c, b, c8, b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, 
        o7, n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, 
        w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, 
        e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, n5, 
        m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, v4, 
        u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4 );
  input h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3,
         p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2,
         y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2,
         h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1,
         q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1,
         z0, y0, x0, w0, v0, u0, t0, s0, r0, o0, n0, m0, l0, k0, j0, i0, h0,
         g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m,
         l, k, j, i, h, g, f, e, d, c, b;
  output c8, b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7,
         l7, k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6,
         u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6,
         d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, n5,
         m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4,
         v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4;
  wire   n1008, n1009, n8, n9, n13, n14, n15, n16, n18, n19, n20, n28, n29,
         n30, n31, n32, n36, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n52, n54, n55, n56, n57, n58, n59, n60, n61, n67, n68,
         n69, n70, n71, n72, n76, n77, n78, n79, n80, n96, n97, n98, n99, n102,
         n103, n104, n105, n106, n112, n113, n114, n115, n118, n119, n120,
         n121, n122, n123, n124, n128, n136, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n186, n188, n189, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n316, n317, n318, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n340, n341,
         n342, n350, n351, n352, n353, n354, n355, n356, n357, n362, n363,
         n364, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n386, n393, n394, n395, n399, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n433, n434, n435, n441, n442, n443,
         n444, n445, n450, n451, n452, n457, n458, n459, n466, n467, n468,
         n469, n470, n471, n476, n477, n478, n479, n480, n485, n487, n488,
         n489, n490, n491, n492, n497, n498, n499, n501, n502, n503, n504,
         n505, n506, n507, n512, n513, n514, n515, n516, n522, n527, n529,
         n530, n531, n532, n533, n534, n535, n536, n541, n542, n543, n544,
         n545, n551, n556, n559, n560, n561, n562, n563, n564, n565, n571,
         n572, n573, n574, n575, n576, n577, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n625, n626, n627, n628, n629, n660, n661, n662,
         n663, n664, n665, n666, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1010, n1011, n1012, n1013, n1014;

  and2 U1 ( .A1(n8), .A2(n9), .Z(z7) );
  and2 U4 ( .A1(n13), .A2(n14), .Z(z6) );
  or2 U5 ( .A1(n15), .A2(n16), .Z(n14) );
  and2 U6 ( .A1(e3), .A2(n712), .Z(n15) );
  and2 U7 ( .A1(n18), .A2(n19), .Z(n13) );
  or2 U8 ( .A1(f3), .A2(n20), .Z(n19) );
  or2 U9 ( .A1(e3), .A2(h), .Z(n18) );
  and2 U15 ( .A1(n28), .A2(n29), .Z(z4) );
  or2 U16 ( .A1(o), .A2(n30), .Z(n29) );
  or2 U17 ( .A1(n31), .A2(n32), .Z(n28) );
  and2 U18 ( .A1(e1), .A2(n1010), .Z(n32) );
  and2 U23 ( .A1(n38), .A2(n39), .Z(y6) );
  or2 U24 ( .A1(n40), .A2(n16), .Z(n39) );
  and2 U25 ( .A1(d3), .A2(n1010), .Z(n40) );
  and2 U26 ( .A1(n41), .A2(n42), .Z(n38) );
  or2 U27 ( .A1(e3), .A2(n20), .Z(n42) );
  or2 U28 ( .A1(d3), .A2(h), .Z(n41) );
  and2 U29 ( .A1(n43), .A2(b), .Z(y5) );
  and2 U30 ( .A1(n44), .A2(n45), .Z(n43) );
  or2 U31 ( .A1(n46), .A2(n1009), .Z(n44) );
  and2 U32 ( .A1(d2), .A2(n1006), .Z(n46) );
  and2 U33 ( .A1(n47), .A2(n48), .Z(y4) );
  or2 U34 ( .A1(n), .A2(n30), .Z(n48) );
  or2 U35 ( .A1(n31), .A2(n49), .Z(n47) );
  and2 U36 ( .A1(d1), .A2(n711), .Z(n49) );
  and2 U37 ( .A1(n50), .A2(n36), .Z(x7) );
  or2 U40 ( .A1(n54), .A2(c4), .Z(n50) );
  and2 U41 ( .A1(n55), .A2(n56), .Z(n54) );
  and2 U42 ( .A1(b4), .A2(a4), .Z(n55) );
  and2 U43 ( .A1(n57), .A2(n58), .Z(x6) );
  or2 U44 ( .A1(n59), .A2(n16), .Z(n58) );
  and2 U45 ( .A1(c3), .A2(n711), .Z(n59) );
  and2 U46 ( .A1(n60), .A2(n61), .Z(n57) );
  or2 U47 ( .A1(d3), .A2(n20), .Z(n61) );
  or2 U48 ( .A1(c3), .A2(h), .Z(n60) );
  and2 U54 ( .A1(n67), .A2(n68), .Z(x4) );
  or2 U55 ( .A1(m), .A2(n30), .Z(n68) );
  or2 U56 ( .A1(n31), .A2(n69), .Z(n67) );
  and2 U57 ( .A1(c1), .A2(n712), .Z(n69) );
  or2 U58 ( .A1(n70), .A2(n71), .Z(w7) );
  and2 U59 ( .A1(b4), .A2(n72), .Z(n71) );
  and2 U63 ( .A1(n76), .A2(n77), .Z(w6) );
  or2 U64 ( .A1(n78), .A2(n16), .Z(n77) );
  and2 U65 ( .A1(b3), .A2(n712), .Z(n78) );
  and2 U66 ( .A1(n79), .A2(n80), .Z(n76) );
  or2 U67 ( .A1(c3), .A2(n20), .Z(n80) );
  or2 U68 ( .A1(b3), .A2(h), .Z(n79) );
  and2 U82 ( .A1(n96), .A2(n97), .Z(w4) );
  or2 U83 ( .A1(l), .A2(n30), .Z(n97) );
  or2 U84 ( .A1(n31), .A2(n98), .Z(n96) );
  and2 U85 ( .A1(b1), .A2(n1010), .Z(n98) );
  and2 U86 ( .A1(n99), .A2(n72), .Z(v7) );
  or2 U89 ( .A1(n56), .A2(a4), .Z(n99) );
  and2 U90 ( .A1(z3), .A2(y3), .Z(n56) );
  and2 U91 ( .A1(n102), .A2(n103), .Z(v6) );
  or2 U92 ( .A1(n104), .A2(n16), .Z(n103) );
  and2 U93 ( .A1(a3), .A2(n1010), .Z(n104) );
  and2 U94 ( .A1(n105), .A2(n106), .Z(n102) );
  or2 U95 ( .A1(b3), .A2(n20), .Z(n106) );
  or2 U96 ( .A1(a3), .A2(h), .Z(n105) );
  and2 U101 ( .A1(n112), .A2(n113), .Z(v4) );
  or2 U102 ( .A1(k), .A2(n30), .Z(n113) );
  or2 U103 ( .A1(n31), .A2(n114), .Z(n112) );
  and2 U104 ( .A1(a1), .A2(n711), .Z(n114) );
  and2 U105 ( .A1(n115), .A2(n52), .Z(u7) );
  or2 U108 ( .A1(y3), .A2(z3), .Z(n115) );
  and2 U109 ( .A1(n118), .A2(n119), .Z(u6) );
  or2 U110 ( .A1(n120), .A2(n16), .Z(n119) );
  and2 U111 ( .A1(z2), .A2(n1010), .Z(n120) );
  and2 U112 ( .A1(n121), .A2(n122), .Z(n118) );
  or2 U113 ( .A1(g), .A2(n123), .Z(n122) );
  or2 U114 ( .A1(z2), .A2(n124), .Z(n121) );
  and2 U122 ( .A1(i2), .A2(r2), .Z(n136) );
  and2 U141 ( .A1(r2), .A2(n165), .Z(n164) );
  and2 U142 ( .A1(n166), .A2(n167), .Z(u4) );
  or2 U143 ( .A1(j), .A2(n30), .Z(n167) );
  or2 U144 ( .A1(n31), .A2(n168), .Z(n166) );
  and2 U145 ( .A1(z0), .A2(n712), .Z(n168) );
  and2 U146 ( .A1(n169), .A2(n170), .Z(t6) );
  or2 U147 ( .A1(n171), .A2(n16), .Z(n170) );
  and2 U148 ( .A1(y2), .A2(n711), .Z(n171) );
  and2 U149 ( .A1(n172), .A2(n173), .Z(n169) );
  or2 U150 ( .A1(z2), .A2(n123), .Z(n173) );
  or2 U151 ( .A1(y2), .A2(n124), .Z(n172) );
  or2 U152 ( .A1(n128), .A2(n0), .Z(t5) );
  and2 U153 ( .A1(n174), .A2(n175), .Z(t4) );
  or2 U154 ( .A1(q), .A2(n176), .Z(n175) );
  or2 U155 ( .A1(n177), .A2(n178), .Z(n174) );
  and2 U156 ( .A1(y0), .A2(n1010), .Z(n178) );
  and2 U157 ( .A1(n179), .A2(n180), .Z(s7) );
  and2 U161 ( .A1(n186), .A2(n1010), .Z(n181) );
  or2 U162 ( .A1(g1), .A2(n708), .Z(n186) );
  and2 U163 ( .A1(n188), .A2(n189), .Z(n179) );
  or2 U164 ( .A1(w1), .A2(n707), .Z(n189) );
  and2 U166 ( .A1(n192), .A2(n193), .Z(s6) );
  or2 U167 ( .A1(n194), .A2(n16), .Z(n193) );
  and2 U168 ( .A1(x2), .A2(n1010), .Z(n194) );
  and2 U169 ( .A1(n195), .A2(n196), .Z(n192) );
  or2 U170 ( .A1(y2), .A2(n123), .Z(n196) );
  or2 U171 ( .A1(x2), .A2(n124), .Z(n195) );
  and2 U172 ( .A1(n197), .A2(n198), .Z(s4) );
  or2 U173 ( .A1(p), .A2(n176), .Z(n198) );
  or2 U174 ( .A1(n177), .A2(n199), .Z(n197) );
  and2 U175 ( .A1(x0), .A2(n712), .Z(n199) );
  and2 U176 ( .A1(n200), .A2(n201), .Z(r7) );
  and2 U182 ( .A1(n208), .A2(n712), .Z(n202) );
  or2 U183 ( .A1(f1), .A2(n708), .Z(n208) );
  and2 U184 ( .A1(n209), .A2(n210), .Z(n200) );
  or2 U185 ( .A1(v1), .A2(n707), .Z(n210) );
  and2 U187 ( .A1(n211), .A2(n212), .Z(r6) );
  or2 U188 ( .A1(n213), .A2(n16), .Z(n212) );
  and2 U189 ( .A1(w2), .A2(n712), .Z(n213) );
  and2 U190 ( .A1(n214), .A2(n215), .Z(n211) );
  or2 U191 ( .A1(x2), .A2(n123), .Z(n215) );
  or2 U192 ( .A1(w2), .A2(n124), .Z(n214) );
  and2 U193 ( .A1(n216), .A2(n217), .Z(r5) );
  or2 U194 ( .A1(a0), .A2(n218), .Z(n217) );
  or2 U195 ( .A1(n219), .A2(n220), .Z(n216) );
  and2 U196 ( .A1(w1), .A2(n1010), .Z(n220) );
  and2 U197 ( .A1(n221), .A2(n222), .Z(r4) );
  or2 U198 ( .A1(o), .A2(n176), .Z(n222) );
  or2 U199 ( .A1(n177), .A2(n223), .Z(n221) );
  and2 U200 ( .A1(w0), .A2(n711), .Z(n223) );
  and2 U201 ( .A1(n224), .A2(n225), .Z(q7) );
  and2 U207 ( .A1(n231), .A2(n1010), .Z(n226) );
  or2 U208 ( .A1(e1), .A2(n708), .Z(n231) );
  and2 U209 ( .A1(n232), .A2(n233), .Z(n224) );
  or2 U210 ( .A1(u1), .A2(n707), .Z(n233) );
  and2 U212 ( .A1(n234), .A2(n235), .Z(q6) );
  or2 U213 ( .A1(n236), .A2(n16), .Z(n235) );
  and2 U214 ( .A1(v2), .A2(n711), .Z(n236) );
  and2 U215 ( .A1(n237), .A2(n238), .Z(n234) );
  or2 U216 ( .A1(w2), .A2(n123), .Z(n238) );
  or2 U217 ( .A1(v2), .A2(n124), .Z(n237) );
  and2 U218 ( .A1(n239), .A2(n240), .Z(q5) );
  or2 U219 ( .A1(z), .A2(n218), .Z(n240) );
  or2 U220 ( .A1(n219), .A2(n241), .Z(n239) );
  and2 U221 ( .A1(v1), .A2(n712), .Z(n241) );
  and2 U222 ( .A1(n242), .A2(n243), .Z(q4) );
  or2 U223 ( .A1(n), .A2(n176), .Z(n243) );
  or2 U224 ( .A1(n177), .A2(n244), .Z(n242) );
  and2 U225 ( .A1(v0), .A2(n1010), .Z(n244) );
  and2 U226 ( .A1(n245), .A2(n246), .Z(p7) );
  and2 U232 ( .A1(n252), .A2(n711), .Z(n247) );
  or2 U233 ( .A1(d1), .A2(n708), .Z(n252) );
  and2 U234 ( .A1(n253), .A2(n254), .Z(n245) );
  or2 U235 ( .A1(t1), .A2(n707), .Z(n254) );
  and2 U237 ( .A1(n255), .A2(n256), .Z(p6) );
  or2 U238 ( .A1(n257), .A2(n16), .Z(n256) );
  and2 U239 ( .A1(u2), .A2(n712), .Z(n257) );
  and2 U240 ( .A1(n258), .A2(n259), .Z(n255) );
  or2 U241 ( .A1(v2), .A2(n123), .Z(n259) );
  or2 U242 ( .A1(u2), .A2(n124), .Z(n258) );
  and2 U243 ( .A1(n260), .A2(n261), .Z(p5) );
  or2 U244 ( .A1(y), .A2(n218), .Z(n261) );
  or2 U245 ( .A1(n219), .A2(n262), .Z(n260) );
  and2 U246 ( .A1(u1), .A2(n711), .Z(n262) );
  and2 U247 ( .A1(n263), .A2(n264), .Z(p4) );
  or2 U248 ( .A1(m), .A2(n176), .Z(n264) );
  or2 U249 ( .A1(n177), .A2(n265), .Z(n263) );
  and2 U250 ( .A1(u0), .A2(n712), .Z(n265) );
  and2 U251 ( .A1(n266), .A2(n267), .Z(o7) );
  and2 U257 ( .A1(n273), .A2(n712), .Z(n268) );
  or2 U258 ( .A1(c1), .A2(n708), .Z(n273) );
  and2 U259 ( .A1(n274), .A2(n275), .Z(n266) );
  or2 U260 ( .A1(s1), .A2(n707), .Z(n275) );
  and2 U262 ( .A1(n276), .A2(n277), .Z(o6) );
  or2 U263 ( .A1(n278), .A2(n16), .Z(n277) );
  and2 U264 ( .A1(t2), .A2(n1010), .Z(n278) );
  and2 U265 ( .A1(n279), .A2(n280), .Z(n276) );
  or2 U266 ( .A1(u2), .A2(n123), .Z(n280) );
  or2 U267 ( .A1(t2), .A2(n124), .Z(n279) );
  and2 U268 ( .A1(n281), .A2(n282), .Z(o5) );
  or2 U269 ( .A1(x), .A2(n218), .Z(n282) );
  or2 U270 ( .A1(n219), .A2(n283), .Z(n281) );
  and2 U271 ( .A1(t1), .A2(n1010), .Z(n283) );
  and2 U272 ( .A1(n284), .A2(n285), .Z(o4) );
  or2 U273 ( .A1(l), .A2(n176), .Z(n285) );
  or2 U274 ( .A1(n177), .A2(n286), .Z(n284) );
  and2 U275 ( .A1(t0), .A2(n1010), .Z(n286) );
  and2 U276 ( .A1(n287), .A2(n288), .Z(n7) );
  and2 U282 ( .A1(n294), .A2(n1010), .Z(n289) );
  or2 U283 ( .A1(b1), .A2(n708), .Z(n294) );
  and2 U284 ( .A1(n295), .A2(n296), .Z(n287) );
  or2 U285 ( .A1(r1), .A2(n707), .Z(n296) );
  and2 U287 ( .A1(n297), .A2(n298), .Z(n6) );
  or2 U288 ( .A1(n299), .A2(n16), .Z(n298) );
  and2 U289 ( .A1(s2), .A2(n712), .Z(n299) );
  and2 U290 ( .A1(n300), .A2(n301), .Z(n297) );
  or2 U291 ( .A1(t2), .A2(n123), .Z(n301) );
  or2 U292 ( .A1(h), .A2(n302), .Z(n123) );
  or2 U293 ( .A1(s2), .A2(n124), .Z(n300) );
  and2 U294 ( .A1(n303), .A2(n304), .Z(n5) );
  or2 U295 ( .A1(w), .A2(n218), .Z(n304) );
  or2 U296 ( .A1(n219), .A2(n305), .Z(n303) );
  and2 U297 ( .A1(s1), .A2(n711), .Z(n305) );
  and2 U298 ( .A1(n306), .A2(n307), .Z(n4) );
  or2 U299 ( .A1(k), .A2(n176), .Z(n307) );
  or2 U300 ( .A1(n177), .A2(n308), .Z(n306) );
  and2 U301 ( .A1(s0), .A2(n711), .Z(n308) );
  and2 U302 ( .A1(n309), .A2(n310), .Z(m7) );
  and2 U308 ( .A1(n316), .A2(n711), .Z(n311) );
  or2 U309 ( .A1(a1), .A2(n708), .Z(n316) );
  and2 U310 ( .A1(n317), .A2(n318), .Z(n309) );
  or2 U311 ( .A1(q1), .A2(n707), .Z(n318) );
  and2 U318 ( .A1(n324), .A2(n325), .Z(m5) );
  or2 U319 ( .A1(v), .A2(n218), .Z(n325) );
  or2 U320 ( .A1(n219), .A2(n326), .Z(n324) );
  and2 U321 ( .A1(r1), .A2(n712), .Z(n326) );
  and2 U322 ( .A1(n327), .A2(n328), .Z(m4) );
  or2 U323 ( .A1(j), .A2(n176), .Z(n328) );
  or2 U324 ( .A1(r), .A2(n329), .Z(n176) );
  or2 U325 ( .A1(n177), .A2(n330), .Z(n327) );
  and2 U326 ( .A1(r0), .A2(n712), .Z(n330) );
  and2 U327 ( .A1(n331), .A2(n332), .Z(n177) );
  and2 U328 ( .A1(n333), .A2(n334), .Z(l7) );
  and2 U334 ( .A1(n340), .A2(n711), .Z(n335) );
  or2 U335 ( .A1(z0), .A2(n708), .Z(n340) );
  and2 U336 ( .A1(n341), .A2(n342), .Z(n333) );
  or2 U337 ( .A1(p1), .A2(n707), .Z(n342) );
  and2 U347 ( .A1(n350), .A2(n351), .Z(l5) );
  or2 U348 ( .A1(u), .A2(n218), .Z(n351) );
  or2 U349 ( .A1(n219), .A2(n352), .Z(n350) );
  and2 U350 ( .A1(q1), .A2(n1010), .Z(n352) );
  and2 U351 ( .A1(n353), .A2(n1006), .Z(l4) );
  or2 U352 ( .A1(n354), .A2(c2), .Z(n353) );
  and2 U353 ( .A1(n355), .A2(n356), .Z(k7) );
  and2 U359 ( .A1(n362), .A2(n712), .Z(n357) );
  or2 U360 ( .A1(y0), .A2(n708), .Z(n362) );
  and2 U361 ( .A1(n363), .A2(n364), .Z(n355) );
  or2 U363 ( .A1(o1), .A2(n707), .Z(n363) );
  and2 U369 ( .A1(n370), .A2(n371), .Z(k5) );
  or2 U370 ( .A1(t), .A2(n218), .Z(n371) );
  or2 U371 ( .A1(n372), .A2(n373), .Z(n218) );
  or2 U372 ( .A1(n219), .A2(n374), .Z(n370) );
  and2 U373 ( .A1(p1), .A2(n711), .Z(n374) );
  and2 U374 ( .A1(b0), .A2(n375), .Z(n219) );
  and2 U376 ( .A1(n378), .A2(n379), .Z(n377) );
  and2 U377 ( .A1(n380), .A2(n381), .Z(n379) );
  and2 U378 ( .A1(n1005), .A2(n711), .Z(n380) );
  or2 U385 ( .A1(r2), .A2(n1007), .Z(n386) );
  or2 U391 ( .A1(q2), .A2(d0), .Z(n393) );
  and2 U395 ( .A1(n394), .A2(n711), .Z(n376) );
  and2 U418 ( .A1(n420), .A2(m0), .Z(n395) );
  and2 U419 ( .A1(a2), .A2(n421), .Z(n420) );
  or2 U420 ( .A1(n422), .A2(n423), .Z(n421) );
  and2 U421 ( .A1(n424), .A2(d0), .Z(n423) );
  and2 U424 ( .A1(n425), .A2(e2), .Z(n422) );
  and2 U425 ( .A1(n165), .A2(n1003), .Z(n425) );
  inv1 U426 ( .I(d0), .ZN(n165) );
  and2 U427 ( .A1(n426), .A2(n427), .Z(j7) );
  and2 U433 ( .A1(n433), .A2(n712), .Z(n428) );
  or2 U434 ( .A1(x0), .A2(n708), .Z(n433) );
  and2 U435 ( .A1(n434), .A2(n435), .Z(n426) );
  or2 U437 ( .A1(n1), .A2(n707), .Z(n434) );
  and2 U443 ( .A1(n441), .A2(n442), .Z(j5) );
  or2 U444 ( .A1(a0), .A2(n443), .Z(n442) );
  or2 U445 ( .A1(n444), .A2(n445), .Z(n441) );
  and2 U446 ( .A1(o1), .A2(n712), .Z(n445) );
  and2 U453 ( .A1(n450), .A2(n451), .Z(i7) );
  and2 U459 ( .A1(n457), .A2(n712), .Z(n452) );
  or2 U460 ( .A1(w0), .A2(n708), .Z(n457) );
  and2 U461 ( .A1(n458), .A2(n459), .Z(n450) );
  or2 U463 ( .A1(m1), .A2(n707), .Z(n458) );
  and2 U471 ( .A1(n466), .A2(n467), .Z(i5) );
  or2 U472 ( .A1(z), .A2(n443), .Z(n467) );
  or2 U473 ( .A1(n444), .A2(n468), .Z(n466) );
  and2 U474 ( .A1(n1), .A2(n712), .Z(n468) );
  inv1 U475 ( .I(n399), .ZN(i4) );
  and2 U476 ( .A1(n381), .A2(x1), .Z(n399) );
  inv1 U477 ( .I(a2), .ZN(n381) );
  and2 U478 ( .A1(n469), .A2(n470), .Z(h7) );
  and2 U484 ( .A1(n476), .A2(n1010), .Z(n471) );
  or2 U485 ( .A1(v0), .A2(n708), .Z(n476) );
  and2 U486 ( .A1(n477), .A2(n478), .Z(n469) );
  or2 U488 ( .A1(l1), .A2(n707), .Z(n477) );
  and2 U489 ( .A1(n479), .A2(n480), .Z(h6) );
  and2 U496 ( .A1(m2), .A2(n711), .Z(n485) );
  and2 U497 ( .A1(n487), .A2(n488), .Z(h5) );
  or2 U498 ( .A1(y), .A2(n443), .Z(n488) );
  or2 U499 ( .A1(n444), .A2(n489), .Z(n487) );
  and2 U500 ( .A1(m1), .A2(n1010), .Z(n489) );
  and2 U501 ( .A1(n490), .A2(n491), .Z(g7) );
  and2 U507 ( .A1(n497), .A2(n711), .Z(n492) );
  or2 U508 ( .A1(u0), .A2(n708), .Z(n497) );
  and2 U509 ( .A1(n498), .A2(n499), .Z(n490) );
  or2 U511 ( .A1(k1), .A2(n707), .Z(n498) );
  and2 U519 ( .A1(l2), .A2(n711), .Z(n501) );
  and2 U520 ( .A1(n502), .A2(n503), .Z(g5) );
  or2 U521 ( .A1(x), .A2(n443), .Z(n503) );
  or2 U522 ( .A1(n444), .A2(n504), .Z(n502) );
  and2 U523 ( .A1(l1), .A2(n1010), .Z(n504) );
  and2 U524 ( .A1(n505), .A2(n506), .Z(f7) );
  and2 U530 ( .A1(n512), .A2(n711), .Z(n507) );
  or2 U531 ( .A1(t0), .A2(n708), .Z(n512) );
  and2 U532 ( .A1(n513), .A2(n514), .Z(n505) );
  or2 U534 ( .A1(j1), .A2(n707), .Z(n513) );
  and2 U535 ( .A1(n515), .A2(n516), .Z(f6) );
  or2 U540 ( .A1(k2), .A2(n1005), .Z(n522) );
  or2 U546 ( .A1(n529), .A2(n530), .Z(n527) );
  and2 U547 ( .A1(n531), .A2(n532), .Z(f5) );
  or2 U548 ( .A1(w), .A2(n443), .Z(n532) );
  or2 U549 ( .A1(n444), .A2(n533), .Z(n531) );
  and2 U550 ( .A1(k1), .A2(n711), .Z(n533) );
  and2 U551 ( .A1(n534), .A2(n535), .Z(e7) );
  and2 U557 ( .A1(n541), .A2(n712), .Z(n536) );
  or2 U558 ( .A1(s0), .A2(n708), .Z(n541) );
  and2 U559 ( .A1(n542), .A2(n543), .Z(n534) );
  or2 U561 ( .A1(i1), .A2(n707), .Z(n542) );
  and2 U562 ( .A1(n544), .A2(n545), .Z(e6) );
  or2 U567 ( .A1(j2), .A2(n1005), .Z(n551) );
  inv1 U573 ( .I(g0), .ZN(n529) );
  inv1 U576 ( .I(n559), .ZN(n556) );
  or2 U577 ( .A1(n530), .A2(o2), .Z(n559) );
  or2 U578 ( .A1(e0), .A2(f0), .Z(n530) );
  and2 U579 ( .A1(n560), .A2(n561), .Z(e5) );
  or2 U580 ( .A1(v), .A2(n443), .Z(n561) );
  or2 U581 ( .A1(n444), .A2(n562), .Z(n560) );
  and2 U582 ( .A1(j1), .A2(n1010), .Z(n562) );
  and2 U583 ( .A1(n563), .A2(n564), .Z(d7) );
  and2 U596 ( .A1(n571), .A2(n1010), .Z(n565) );
  or2 U597 ( .A1(r0), .A2(n708), .Z(n571) );
  and2 U599 ( .A1(n1014), .A2(d), .Z(n572) );
  and2 U600 ( .A1(n573), .A2(n574), .Z(n563) );
  inv1 U603 ( .I(c), .ZN(n575) );
  or2 U605 ( .A1(h1), .A2(n707), .Z(n573) );
  inv1 U607 ( .I(n576), .ZN(d6) );
  or2 U608 ( .A1(n577), .A2(y1), .Z(n576) );
  and2 U626 ( .A1(n585), .A2(n586), .Z(d5) );
  or2 U627 ( .A1(u), .A2(n443), .Z(n586) );
  or2 U628 ( .A1(n444), .A2(n587), .Z(n585) );
  and2 U629 ( .A1(i1), .A2(n712), .Z(n587) );
  and2 U630 ( .A1(n588), .A2(n589), .Z(c8) );
  and2 U631 ( .A1(n45), .A2(n1006), .Z(n589) );
  inv1 U632 ( .I(n354), .ZN(n45) );
  and2 U633 ( .A1(g2), .A2(h2), .Z(n354) );
  and2 U634 ( .A1(b), .A2(n590), .Z(n588) );
  or2 U635 ( .A1(n591), .A2(h4), .Z(n590) );
  and2 U636 ( .A1(l0), .A2(d2), .Z(n591) );
  and2 U637 ( .A1(n592), .A2(n593), .Z(c7) );
  or2 U638 ( .A1(n594), .A2(n16), .Z(n593) );
  and2 U639 ( .A1(h3), .A2(n711), .Z(n594) );
  and2 U640 ( .A1(n595), .A2(n596), .Z(n592) );
  or2 U641 ( .A1(g), .A2(n20), .Z(n596) );
  or2 U642 ( .A1(h), .A2(h3), .Z(n595) );
  and2 U643 ( .A1(n1006), .A2(l0), .Z(n1009) );
  and2 U644 ( .A1(n597), .A2(n598), .Z(c5) );
  or2 U645 ( .A1(t), .A2(n443), .Z(n598) );
  or2 U646 ( .A1(b0), .A2(n373), .Z(n443) );
  inv1 U647 ( .I(s), .ZN(n373) );
  or2 U648 ( .A1(n444), .A2(n599), .Z(n597) );
  and2 U649 ( .A1(h1), .A2(n711), .Z(n599) );
  and2 U650 ( .A1(n372), .A2(n375), .Z(n444) );
  and2 U651 ( .A1(n712), .A2(s), .Z(n375) );
  inv1 U652 ( .I(b0), .ZN(n372) );
  and2 U653 ( .A1(n1002), .A2(n600), .Z(b8) );
  or2 U654 ( .A1(n601), .A2(n602), .Z(n600) );
  inv1 U655 ( .I(n603), .ZN(n602) );
  or2 U656 ( .A1(n604), .A2(g4), .Z(n603) );
  and2 U657 ( .A1(g4), .A2(n604), .Z(n601) );
  and2 U660 ( .A1(n608), .A2(n609), .Z(b7) );
  or2 U661 ( .A1(n610), .A2(n16), .Z(n609) );
  and2 U662 ( .A1(g3), .A2(n711), .Z(n610) );
  and2 U663 ( .A1(n611), .A2(n612), .Z(n608) );
  or2 U664 ( .A1(h3), .A2(n20), .Z(n612) );
  or2 U665 ( .A1(g3), .A2(h), .Z(n611) );
  and2 U666 ( .A1(h2), .A2(n1006), .Z(b6) );
  and2 U667 ( .A1(n613), .A2(n614), .Z(b5) );
  or2 U668 ( .A1(q), .A2(n30), .Z(n614) );
  or2 U669 ( .A1(n31), .A2(n615), .Z(n613) );
  and2 U670 ( .A1(g1), .A2(n711), .Z(n615) );
  and2 U671 ( .A1(n616), .A2(n617), .Z(a8) );
  and2 U685 ( .A1(n625), .A2(n626), .Z(a7) );
  or2 U686 ( .A1(n627), .A2(n16), .Z(n626) );
  and2 U687 ( .A1(n1010), .A2(f), .Z(n16) );
  and2 U688 ( .A1(f3), .A2(n1010), .Z(n627) );
  and2 U689 ( .A1(n628), .A2(n629), .Z(n625) );
  or2 U690 ( .A1(g3), .A2(n20), .Z(n629) );
  or2 U691 ( .A1(n302), .A2(n124), .Z(n20) );
  inv1 U692 ( .I(h), .ZN(n124) );
  inv1 U693 ( .I(f), .ZN(n302) );
  or2 U694 ( .A1(f3), .A2(h), .Z(n628) );
  and2 U745 ( .A1(n660), .A2(n661), .Z(a5) );
  or2 U746 ( .A1(p), .A2(n30), .Z(n661) );
  or2 U747 ( .A1(n329), .A2(n331), .Z(n30) );
  inv1 U748 ( .I(r), .ZN(n331) );
  inv1 U749 ( .I(i), .ZN(n329) );
  or2 U750 ( .A1(n31), .A2(n662), .Z(n660) );
  and2 U751 ( .A1(f1), .A2(n712), .Z(n662) );
  and2 U752 ( .A1(r), .A2(n332), .Z(n31) );
  and2 U753 ( .A1(n711), .A2(i), .Z(n332) );
  and2 U757 ( .A1(n665), .A2(a2), .Z(n664) );
  inv1 U758 ( .I(n923), .ZN(n665) );
  buf0 U761 ( .I(n1009), .Z(c6) );
  buf0 U762 ( .I(n1008), .Z(t7) );
  inv1 U764 ( .I(n669), .ZN(n781) );
  or2 U766 ( .A1(n982), .A2(n673), .Z(n671) );
  and2 U767 ( .A1(n671), .A2(n672), .Z(n989) );
  or2 U768 ( .A1(r2), .A2(n690), .Z(n672) );
  or2 U769 ( .A1(i2), .A2(r2), .Z(n673) );
  and2 U770 ( .A1(n971), .A2(o2), .Z(n674) );
  and2 U771 ( .A1(o2), .A2(n966), .Z(n675) );
  and2 U775 ( .A1(n677), .A2(n678), .Z(n881) );
  or2 U776 ( .A1(n128), .A2(n880), .Z(n678) );
  or2 U777 ( .A1(n884), .A2(n128), .Z(n679) );
  inv1 U779 ( .I(n884), .ZN(n681) );
  or2 U782 ( .A1(n959), .A2(f2), .Z(n684) );
  and2 U788 ( .A1(n985), .A2(n690), .Z(n689) );
  inv1 U790 ( .I(n984), .ZN(n690) );
  or2 U791 ( .A1(n898), .A2(n693), .Z(n691) );
  or2 U793 ( .A1(z1), .A2(n1005), .Z(n692) );
  or2 U794 ( .A1(n897), .A2(z1), .Z(n693) );
  and2 U796 ( .A1(n675), .A2(n967), .Z(n695) );
  inv1 U797 ( .I(n674), .ZN(n978) );
  inv1 U805 ( .I(n953), .ZN(n702) );
  inv1 U808 ( .I(n865), .ZN(n705) );
  inv1 U809 ( .I(n705), .ZN(n706) );
  inv1 U810 ( .I(e), .ZN(n707) );
  inv1 U811 ( .I(n572), .ZN(n708) );
  inv1 U814 ( .I(y1), .ZN(n711) );
  inv1 U815 ( .I(y1), .ZN(n712) );
  inv1 U816 ( .I(y3), .ZN(n713) );
  inv1 U817 ( .I(f4), .ZN(n939) );
  or2 U818 ( .A1(n713), .A2(n939), .Z(n718) );
  inv1 U819 ( .I(b4), .ZN(n851) );
  inv1 U820 ( .I(c4), .ZN(n714) );
  or2 U821 ( .A1(n851), .A2(n714), .Z(n854) );
  inv1 U822 ( .I(z3), .ZN(n859) );
  or2 U823 ( .A1(n854), .A2(n859), .Z(n717) );
  or2 U825 ( .A1(d4), .A2(n938), .Z(n715) );
  inv1 U826 ( .I(a4), .ZN(n860) );
  or2 U827 ( .A1(n715), .A2(n860), .Z(n716) );
  or2 U828 ( .A1(n717), .A2(n716), .Z(n863) );
  or2 U829 ( .A1(n718), .A2(n863), .Z(n604) );
  inv1 U831 ( .I(n994), .ZN(n1002) );
  and2 U832 ( .A1(n604), .A2(n1002), .Z(n616) );
  inv1 U833 ( .I(n863), .ZN(n719) );
  and2 U834 ( .A1(y3), .A2(n719), .Z(n720) );
  or2 U835 ( .A1(n720), .A2(f4), .Z(n617) );
  inv1 U836 ( .I(n0), .ZN(n1006) );
  inv1 U838 ( .I(p2), .ZN(n977) );
  and2 U839 ( .A1(g0), .A2(n977), .Z(n721) );
  or2 U840 ( .A1(n721), .A2(o2), .Z(n723) );
  inv1 U841 ( .I(o2), .ZN(n973) );
  or2 U842 ( .A1(n973), .A2(p2), .Z(n722) );
  inv1 U844 ( .I(j2), .ZN(n739) );
  and2 U845 ( .A1(o2), .A2(n739), .Z(n725) );
  inv1 U847 ( .I(n2), .ZN(n787) );
  or2 U852 ( .A1(n981), .A2(x1), .Z(n727) );
  and2 U853 ( .A1(n804), .A2(n727), .Z(n577) );
  or2 U854 ( .A1(e), .A2(d), .Z(n730) );
  or2 U855 ( .A1(n730), .A2(n575), .Z(n840) );
  or2 U856 ( .A1(n840), .A2(s2), .Z(n574) );
  or2 U860 ( .A1(n703), .A2(j3), .Z(n729) );
  or2 U861 ( .A1(n1013), .A2(i3), .Z(n728) );
  and2 U862 ( .A1(n729), .A2(n728), .Z(n731) );
  or2 U863 ( .A1(n730), .A2(c), .Z(n865) );
  or2 U864 ( .A1(n731), .A2(n706), .Z(n732) );
  and2 U865 ( .A1(n565), .A2(n732), .Z(n564) );
  inv1 U866 ( .I(x1), .ZN(n1005) );
  and2 U867 ( .A1(n529), .A2(n973), .Z(n733) );
  or2 U868 ( .A1(n733), .A2(n556), .Z(n736) );
  or2 U869 ( .A1(n734), .A2(p2), .Z(n735) );
  or2 U870 ( .A1(n736), .A2(n735), .Z(n740) );
  inv1 U871 ( .I(n740), .ZN(n737) );
  or2 U872 ( .A1(n737), .A2(j2), .Z(n738) );
  and2 U873 ( .A1(n551), .A2(n738), .Z(n544) );
  or2 U874 ( .A1(x1), .A2(n739), .Z(n741) );
  or2 U875 ( .A1(n741), .A2(n740), .Z(n742) );
  and2 U876 ( .A1(n711), .A2(n742), .Z(n545) );
  or2 U877 ( .A1(n840), .A2(t2), .Z(n543) );
  or2 U878 ( .A1(n703), .A2(k3), .Z(n744) );
  or2 U879 ( .A1(n1012), .A2(j3), .Z(n743) );
  and2 U880 ( .A1(n744), .A2(n743), .Z(n745) );
  or2 U881 ( .A1(n745), .A2(n706), .Z(n746) );
  and2 U882 ( .A1(n536), .A2(n746), .Z(n535) );
  and2 U883 ( .A1(n527), .A2(n977), .Z(n749) );
  or2 U884 ( .A1(n747), .A2(o2), .Z(n748) );
  or2 U885 ( .A1(n749), .A2(n748), .Z(n753) );
  inv1 U886 ( .I(n753), .ZN(n750) );
  or2 U887 ( .A1(n750), .A2(k2), .Z(n751) );
  and2 U888 ( .A1(n522), .A2(n751), .Z(n515) );
  inv1 U889 ( .I(k2), .ZN(n752) );
  or2 U890 ( .A1(x1), .A2(n752), .Z(n754) );
  or2 U891 ( .A1(n754), .A2(n753), .Z(n755) );
  and2 U892 ( .A1(n712), .A2(n755), .Z(n516) );
  or2 U893 ( .A1(n840), .A2(u2), .Z(n514) );
  or2 U894 ( .A1(n704), .A2(l3), .Z(n757) );
  or2 U895 ( .A1(n1012), .A2(k3), .Z(n756) );
  and2 U896 ( .A1(n757), .A2(n756), .Z(n758) );
  or2 U897 ( .A1(n758), .A2(n706), .Z(n759) );
  and2 U898 ( .A1(n507), .A2(n759), .Z(n506) );
  or2 U899 ( .A1(n840), .A2(v2), .Z(n499) );
  or2 U900 ( .A1(n703), .A2(m3), .Z(n761) );
  or2 U901 ( .A1(n1012), .A2(l3), .Z(n760) );
  and2 U902 ( .A1(n761), .A2(n760), .Z(n762) );
  or2 U903 ( .A1(n762), .A2(n706), .Z(n763) );
  and2 U904 ( .A1(n492), .A2(n763), .Z(n491) );
  and2 U906 ( .A1(n712), .A2(n962), .Z(n963) );
  inv1 U907 ( .I(n963), .ZN(s5) );
  or2 U908 ( .A1(n963), .A2(n485), .Z(n479) );
  and2 U909 ( .A1(m2), .A2(n962), .Z(n764) );
  or2 U910 ( .A1(n764), .A2(n788), .Z(n766) );
  inv1 U911 ( .I(m2), .ZN(n782) );
  or2 U912 ( .A1(l2), .A2(n782), .Z(n765) );
  and2 U913 ( .A1(n766), .A2(n765), .Z(n767) );
  inv1 U914 ( .I(n767), .ZN(n480) );
  or2 U915 ( .A1(n840), .A2(w2), .Z(n478) );
  or2 U916 ( .A1(n703), .A2(n3), .Z(n769) );
  or2 U917 ( .A1(n687), .A2(m3), .Z(n768) );
  and2 U918 ( .A1(n769), .A2(n768), .Z(n770) );
  or2 U919 ( .A1(n770), .A2(n706), .Z(n771) );
  and2 U920 ( .A1(n471), .A2(n771), .Z(n470) );
  or2 U921 ( .A1(n840), .A2(x2), .Z(n459) );
  or2 U922 ( .A1(n704), .A2(o3), .Z(n773) );
  or2 U923 ( .A1(n1013), .A2(n3), .Z(n772) );
  and2 U924 ( .A1(n773), .A2(n772), .Z(n774) );
  or2 U925 ( .A1(n774), .A2(n706), .Z(n775) );
  and2 U926 ( .A1(n452), .A2(n775), .Z(n451) );
  or2 U927 ( .A1(n840), .A2(y2), .Z(n435) );
  or2 U928 ( .A1(n704), .A2(p3), .Z(n777) );
  or2 U929 ( .A1(n1013), .A2(o3), .Z(n776) );
  and2 U930 ( .A1(n777), .A2(n776), .Z(n778) );
  or2 U931 ( .A1(n778), .A2(n706), .Z(n779) );
  and2 U932 ( .A1(n428), .A2(n779), .Z(n427) );
  inv1 U933 ( .I(f2), .ZN(n1003) );
  inv1 U934 ( .I(e2), .ZN(n1004) );
  inv1 U935 ( .I(q2), .ZN(n983) );
  inv1 U936 ( .I(r2), .ZN(n990) );
  or2 U940 ( .A1(n399), .A2(n781), .Z(n795) );
  and2 U941 ( .A1(n782), .A2(n2), .Z(n786) );
  and2 U942 ( .A1(h0), .A2(l2), .Z(n784) );
  or2 U944 ( .A1(n784), .A2(n783), .Z(n785) );
  and2 U945 ( .A1(n786), .A2(n785), .Z(n793) );
  and2 U946 ( .A1(m2), .A2(n787), .Z(n791) );
  and2 U947 ( .A1(j0), .A2(l2), .Z(n789) );
  or2 U948 ( .A1(n789), .A2(n682), .Z(n790) );
  and2 U949 ( .A1(n791), .A2(n790), .Z(n792) );
  or2 U952 ( .A1(o2), .A2(p2), .Z(n884) );
  inv1 U955 ( .I(c0), .ZN(n1007) );
  and2 U956 ( .A1(r2), .A2(i2), .Z(n798) );
  inv1 U957 ( .I(i3), .ZN(n797) );
  or2 U958 ( .A1(n798), .A2(n797), .Z(n799) );
  inv1 U959 ( .I(n799), .ZN(n801) );
  and2 U960 ( .A1(n393), .A2(n871), .Z(n800) );
  or2 U961 ( .A1(n801), .A2(n800), .Z(n802) );
  and2 U962 ( .A1(n879), .A2(n802), .Z(n807) );
  inv1 U963 ( .I(z1), .ZN(n874) );
  or2 U964 ( .A1(n990), .A2(n874), .Z(n803) );
  and2 U965 ( .A1(n386), .A2(n803), .Z(n805) );
  or2 U967 ( .A1(n805), .A2(n868), .Z(n806) );
  and2 U968 ( .A1(n807), .A2(n806), .Z(n378) );
  or2 U969 ( .A1(n840), .A2(z2), .Z(n364) );
  or2 U970 ( .A1(n704), .A2(q3), .Z(n809) );
  or2 U971 ( .A1(n1012), .A2(p3), .Z(n808) );
  and2 U972 ( .A1(n809), .A2(n808), .Z(n810) );
  or2 U973 ( .A1(n810), .A2(n706), .Z(n811) );
  and2 U974 ( .A1(n357), .A2(n811), .Z(n356) );
  or2 U975 ( .A1(n840), .A2(a3), .Z(n341) );
  or2 U976 ( .A1(n704), .A2(r3), .Z(n813) );
  or2 U977 ( .A1(n1013), .A2(q3), .Z(n812) );
  and2 U978 ( .A1(n813), .A2(n812), .Z(n814) );
  or2 U979 ( .A1(n814), .A2(n706), .Z(n815) );
  and2 U980 ( .A1(n335), .A2(n815), .Z(n334) );
  or2 U981 ( .A1(n840), .A2(b3), .Z(n317) );
  or2 U982 ( .A1(n704), .A2(s3), .Z(n817) );
  or2 U983 ( .A1(n1012), .A2(r3), .Z(n816) );
  and2 U984 ( .A1(n817), .A2(n816), .Z(n818) );
  or2 U985 ( .A1(n818), .A2(n706), .Z(n819) );
  and2 U986 ( .A1(n311), .A2(n819), .Z(n310) );
  or2 U987 ( .A1(n840), .A2(c3), .Z(n295) );
  or2 U988 ( .A1(n703), .A2(t3), .Z(n821) );
  or2 U989 ( .A1(n687), .A2(s3), .Z(n820) );
  and2 U990 ( .A1(n821), .A2(n820), .Z(n822) );
  or2 U991 ( .A1(n822), .A2(n706), .Z(n823) );
  and2 U992 ( .A1(n289), .A2(n823), .Z(n288) );
  or2 U993 ( .A1(n840), .A2(d3), .Z(n274) );
  or2 U994 ( .A1(n704), .A2(u3), .Z(n825) );
  or2 U995 ( .A1(n1013), .A2(t3), .Z(n824) );
  and2 U996 ( .A1(n825), .A2(n824), .Z(n826) );
  or2 U997 ( .A1(n826), .A2(n706), .Z(n827) );
  and2 U998 ( .A1(n268), .A2(n827), .Z(n267) );
  or2 U999 ( .A1(n840), .A2(e3), .Z(n253) );
  or2 U1000 ( .A1(n704), .A2(v3), .Z(n829) );
  or2 U1001 ( .A1(n1012), .A2(u3), .Z(n828) );
  and2 U1002 ( .A1(n829), .A2(n828), .Z(n830) );
  or2 U1003 ( .A1(n830), .A2(n706), .Z(n831) );
  and2 U1004 ( .A1(n247), .A2(n831), .Z(n246) );
  or2 U1005 ( .A1(n840), .A2(f3), .Z(n232) );
  or2 U1006 ( .A1(n703), .A2(w3), .Z(n833) );
  or2 U1007 ( .A1(n1012), .A2(v3), .Z(n832) );
  and2 U1008 ( .A1(n833), .A2(n832), .Z(n834) );
  and2 U1010 ( .A1(n226), .A2(n835), .Z(n225) );
  or2 U1011 ( .A1(n840), .A2(g3), .Z(n209) );
  or2 U1012 ( .A1(n703), .A2(x3), .Z(n837) );
  or2 U1013 ( .A1(n1013), .A2(w3), .Z(n836) );
  and2 U1014 ( .A1(n837), .A2(n836), .Z(n838) );
  and2 U1016 ( .A1(n202), .A2(n839), .Z(n201) );
  or2 U1017 ( .A1(n840), .A2(h3), .Z(n188) );
  and2 U1018 ( .A1(x3), .A2(n703), .Z(n842) );
  or2 U1019 ( .A1(n842), .A2(n706), .Z(n843) );
  and2 U1020 ( .A1(n181), .A2(n843), .Z(n180) );
  or2 U1021 ( .A1(x1), .A2(n990), .Z(n844) );
  inv1 U1023 ( .I(n845), .ZN(n128) );
  or2 U1024 ( .A1(n994), .A2(y3), .Z(n846) );
  inv1 U1025 ( .I(n846), .ZN(n1008) );
  or2 U1026 ( .A1(n994), .A2(z3), .Z(n847) );
  inv1 U1027 ( .I(n847), .ZN(n848) );
  or2 U1028 ( .A1(n1008), .A2(n848), .Z(n52) );
  or2 U1030 ( .A1(n994), .A2(a4), .Z(n849) );
  inv1 U1032 ( .I(n857), .ZN(n72) );
  and2 U1033 ( .A1(n56), .A2(a4), .Z(n853) );
  and2 U1034 ( .A1(n851), .A2(n1002), .Z(n852) );
  and2 U1035 ( .A1(n853), .A2(n852), .Z(n70) );
  inv1 U1036 ( .I(n854), .ZN(n855) );
  or2 U1037 ( .A1(n994), .A2(n855), .Z(n856) );
  inv1 U1039 ( .I(n997), .ZN(n36) );
  or2 U1042 ( .A1(n860), .A2(n859), .Z(n861) );
  inv1 U1044 ( .I(n996), .ZN(n936) );
  and2 U1045 ( .A1(n998), .A2(n936), .Z(n862) );
  or2 U1046 ( .A1(n862), .A2(e4), .Z(n8) );
  and2 U1047 ( .A1(n863), .A2(n1002), .Z(n864) );
  or2 U1048 ( .A1(n864), .A2(n1008), .Z(n9) );
  or2 U1049 ( .A1(n128), .A2(o0), .Z(n866) );
  and2 U1050 ( .A1(n705), .A2(n866), .Z(n867) );
  or2 U1051 ( .A1(n867), .A2(y1), .Z(j4) );
  and2 U1052 ( .A1(n164), .A2(i2), .Z(n870) );
  inv1 U1053 ( .I(n868), .ZN(n889) );
  and2 U1054 ( .A1(c0), .A2(n889), .Z(n869) );
  or2 U1055 ( .A1(n870), .A2(n869), .Z(n878) );
  or2 U1056 ( .A1(n871), .A2(n885), .Z(n872) );
  or2 U1057 ( .A1(n872), .A2(i3), .Z(n873) );
  inv1 U1058 ( .I(n873), .ZN(n876) );
  or2 U1059 ( .A1(x1), .A2(n874), .Z(n875) );
  or2 U1060 ( .A1(n876), .A2(n875), .Z(n877) );
  or2 U1061 ( .A1(n878), .A2(n877), .Z(n882) );
  inv1 U1062 ( .I(n879), .ZN(n880) );
  and2 U1065 ( .A1(n885), .A2(n892), .Z(n886) );
  and2 U1066 ( .A1(n681), .A2(n886), .Z(n887) );
  and2 U1067 ( .A1(n888), .A2(n887), .Z(n898) );
  and2 U1068 ( .A1(d0), .A2(n136), .Z(n896) );
  and2 U1069 ( .A1(n1007), .A2(n889), .Z(n894) );
  or2 U1073 ( .A1(n896), .A2(n895), .Z(n897) );
  inv1 U1076 ( .I(j0), .ZN(n902) );
  and2 U1077 ( .A1(n902), .A2(f4), .Z(n907) );
  inv1 U1079 ( .I(k0), .ZN(n903) );
  and2 U1080 ( .A1(g4), .A2(n903), .Z(n904) );
  inv1 U1083 ( .I(g4), .ZN(n940) );
  and2 U1084 ( .A1(n940), .A2(k0), .Z(n910) );
  inv1 U1085 ( .I(i0), .ZN(n908) );
  and2 U1086 ( .A1(n908), .A2(e4), .Z(n909) );
  or2 U1087 ( .A1(n910), .A2(n909), .Z(n914) );
  inv1 U1089 ( .I(h4), .ZN(n911) );
  or2 U1090 ( .A1(n912), .A2(n911), .Z(n913) );
  inv1 U1093 ( .I(h0), .ZN(n917) );
  or2 U1094 ( .A1(d4), .A2(n917), .Z(n919) );
  and2 U1096 ( .A1(n919), .A2(n918), .Z(n920) );
  inv1 U1098 ( .I(n922), .ZN(n954) );
  and2 U1099 ( .A1(e2), .A2(f2), .Z(n923) );
  or2 U1100 ( .A1(j0), .A2(i0), .Z(n924) );
  or2 U1101 ( .A1(n924), .A2(k0), .Z(n927) );
  or2 U1105 ( .A1(n664), .A2(n952), .Z(n929) );
  or2 U1106 ( .A1(n954), .A2(n929), .Z(n930) );
  and2 U1107 ( .A1(n1010), .A2(n930), .Z(v5) );
  inv1 U1108 ( .I(b2), .ZN(n931) );
  or2 U1109 ( .A1(n931), .A2(n998), .Z(n932) );
  or2 U1110 ( .A1(n996), .A2(n932), .Z(n935) );
  or2 U1111 ( .A1(f4), .A2(e4), .Z(n933) );
  or2 U1112 ( .A1(g4), .A2(n933), .Z(n934) );
  or2 U1113 ( .A1(n935), .A2(n934), .Z(n949) );
  and2 U1114 ( .A1(n1002), .A2(n949), .Z(n945) );
  and2 U1115 ( .A1(d4), .A2(n936), .Z(n937) );
  and2 U1117 ( .A1(n940), .A2(n939), .Z(n941) );
  and2 U1118 ( .A1(n942), .A2(n941), .Z(n943) );
  or2 U1119 ( .A1(n943), .A2(b2), .Z(n944) );
  and2 U1120 ( .A1(n945), .A2(n944), .Z(w5) );
  inv1 U1121 ( .I(n949), .ZN(n946) );
  or2 U1122 ( .A1(n946), .A2(c2), .Z(n947) );
  and2 U1123 ( .A1(n1002), .A2(n947), .Z(n951) );
  inv1 U1124 ( .I(c2), .ZN(n948) );
  or2 U1125 ( .A1(n949), .A2(n948), .Z(n950) );
  and2 U1126 ( .A1(n951), .A2(n950), .Z(x5) );
  or2 U1127 ( .A1(a2), .A2(n952), .Z(n953) );
  and2 U1128 ( .A1(e2), .A2(n701), .Z(n957) );
  and2 U1131 ( .A1(n1006), .A2(n958), .Z(z5) );
  inv1 U1132 ( .I(n686), .ZN(n959) );
  or2 U1133 ( .A1(n960), .A2(n1003), .Z(n961) );
  inv1 U1135 ( .I(n967), .ZN(n965) );
  or2 U1136 ( .A1(n963), .A2(n501), .Z(n964) );
  and2 U1137 ( .A1(n965), .A2(n964), .Z(g6) );
  and2 U1138 ( .A1(m2), .A2(n2), .Z(n966) );
  inv1 U1140 ( .I(n971), .ZN(n974) );
  and2 U1141 ( .A1(n1010), .A2(n974), .Z(n970) );
  and2 U1142 ( .A1(m2), .A2(n967), .Z(n968) );
  or2 U1143 ( .A1(n968), .A2(n2), .Z(n969) );
  and2 U1144 ( .A1(n970), .A2(n969), .Z(i6) );
  or2 U1145 ( .A1(n971), .A2(o2), .Z(n972) );
  and2 U1146 ( .A1(n711), .A2(n972), .Z(n975) );
  and2 U1147 ( .A1(n975), .A2(n978), .Z(j6) );
  or2 U1148 ( .A1(n695), .A2(p2), .Z(n976) );
  and2 U1149 ( .A1(n712), .A2(n976), .Z(n980) );
  or2 U1150 ( .A1(n978), .A2(n977), .Z(n979) );
  and2 U1151 ( .A1(n980), .A2(n979), .Z(k6) );
  inv1 U1152 ( .I(n981), .ZN(n982) );
  or2 U1154 ( .A1(x1), .A2(n983), .Z(n984) );
  and2 U1155 ( .A1(n712), .A2(n991), .Z(n988) );
  and2 U1156 ( .A1(n1005), .A2(n985), .Z(n986) );
  or2 U1157 ( .A1(n986), .A2(q2), .Z(n987) );
  and2 U1159 ( .A1(n1010), .A2(n989), .Z(n993) );
  or2 U1160 ( .A1(n991), .A2(n990), .Z(n992) );
  and2 U1161 ( .A1(n993), .A2(n992), .Z(m6) );
  or2 U1162 ( .A1(d4), .A2(n994), .Z(n995) );
  or2 U1163 ( .A1(n996), .A2(n995), .Z(n1000) );
  or2 U1164 ( .A1(n998), .A2(n997), .Z(n999) );
  and2 U1165 ( .A1(n1000), .A2(n999), .Z(n1001) );
  inv1 U1166 ( .I(n1001), .ZN(y7) );
  inv1f U755 ( .I(l2), .ZN(n788) );
  or2f U756 ( .A1(n794), .A2(n679), .Z(n677) );
  inv1 U759 ( .I(n694), .ZN(n871) );
  and2 U760 ( .A1(n696), .A2(n697), .Z(n686) );
  and2 U763 ( .A1(n857), .A2(n856), .Z(n997) );
  or2f U765 ( .A1(n376), .A2(n377), .Z(k4) );
  inv1f U772 ( .I(n928), .ZN(n952) );
  and2f U773 ( .A1(n1004), .A2(n955), .Z(n956) );
  or2f U774 ( .A1(n907), .A2(n906), .Z(n916) );
  or2f U778 ( .A1(n0), .A2(l0), .Z(n994) );
  and2f U780 ( .A1(n850), .A2(n849), .Z(n857) );
  inv1f U781 ( .I(n52), .ZN(n850) );
  and2 U783 ( .A1(i0), .A2(n938), .Z(n912) );
  or2 U784 ( .A1(n879), .A2(a2), .Z(n669) );
  inv1 U785 ( .I(n888), .ZN(n794) );
  or2 U786 ( .A1(n780), .A2(n804), .Z(n892) );
  or2 U787 ( .A1(n925), .A2(h0), .Z(n926) );
  inv1 U789 ( .I(n701), .ZN(n955) );
  inv1 U792 ( .I(n689), .ZN(n991) );
  or2 U795 ( .A1(n834), .A2(n706), .Z(n835) );
  or2 U798 ( .A1(n838), .A2(n706), .Z(n839) );
  inv1 U799 ( .I(d4), .ZN(n998) );
  and2 U800 ( .A1(n684), .A2(n685), .Z(a6) );
  inv1 U801 ( .I(y1), .ZN(n1010) );
  or2f U802 ( .A1(n998), .A2(h0), .Z(n918) );
  inv1f U803 ( .I(n688), .ZN(n1011) );
  inv1f U804 ( .I(n1011), .ZN(n1012) );
  inv1f U806 ( .I(n1011), .ZN(n1013) );
  and2f U807 ( .A1(n938), .A2(n937), .Z(n942) );
  inv1 U812 ( .I(n663), .ZN(n700) );
  inv1f U813 ( .I(n841), .ZN(n687) );
  and2 U824 ( .A1(i3), .A2(n890), .Z(n891) );
  or2f U830 ( .A1(n871), .A2(n890), .Z(n879) );
  or2f U837 ( .A1(n724), .A2(m2), .Z(n747) );
  inv1f U843 ( .I(i2), .ZN(n804) );
  and2f U846 ( .A1(f2), .A2(n1004), .Z(n424) );
  or2 U848 ( .A1(n916), .A2(n1004), .Z(n670) );
  and2f U849 ( .A1(n961), .A2(n1006), .Z(n685) );
  or2f U850 ( .A1(n905), .A2(n904), .Z(n906) );
  and2f U851 ( .A1(j0), .A2(n939), .Z(n905) );
  or2f U857 ( .A1(n1004), .A2(n702), .Z(n697) );
  or2f U858 ( .A1(n395), .A2(n796), .Z(n394) );
  and2f U859 ( .A1(n795), .A2(n680), .Z(n796) );
  or2f U905 ( .A1(n700), .A2(n699), .Z(n683) );
  or2f U937 ( .A1(n861), .A2(n920), .Z(n699) );
  and2f U938 ( .A1(n901), .A2(n900), .Z(u5) );
  and2f U939 ( .A1(n711), .A2(n883), .Z(n901) );
  or2f U943 ( .A1(n882), .A2(n881), .Z(n883) );
  or2f U950 ( .A1(n982), .A2(i2), .Z(n985) );
  or2f U951 ( .A1(n726), .A2(n734), .Z(n981) );
  and2f U953 ( .A1(n723), .A2(n722), .Z(n726) );
  or2f U954 ( .A1(n725), .A2(n747), .Z(n734) );
  inv1 U966 ( .I(e), .ZN(n1014) );
  and2f U1009 ( .A1(n967), .A2(n966), .Z(n971) );
  and2f U1015 ( .A1(l2), .A2(n962), .Z(n967) );
  or2f U1022 ( .A1(n865), .A2(n1005), .Z(n962) );
  or2f U1029 ( .A1(n899), .A2(n128), .Z(n900) );
  and2f U1031 ( .A1(n691), .A2(n692), .Z(n899) );
  inv1f U1038 ( .I(n890), .ZN(n885) );
  or2f U1040 ( .A1(j2), .A2(k2), .Z(n890) );
  and2f U1041 ( .A1(n988), .A2(n987), .Z(l6) );
  and2f U1043 ( .A1(n858), .A2(y3), .Z(n663) );
  and2f U1063 ( .A1(c4), .A2(b4), .Z(n858) );
  or2f U1064 ( .A1(n700), .A2(n861), .Z(n996) );
  or2f U1070 ( .A1(n683), .A2(n698), .Z(n696) );
  or2f U1071 ( .A1(n916), .A2(n915), .Z(n921) );
  inv1f U1072 ( .I(n687), .ZN(n703) );
  inv1f U1074 ( .I(n841), .ZN(n688) );
  or2f U1075 ( .A1(n844), .A2(n868), .Z(n845) );
  or2f U1078 ( .A1(n804), .A2(n983), .Z(n868) );
  inv1f U1081 ( .I(n676), .ZN(n780) );
  or2f U1082 ( .A1(q2), .A2(r2), .Z(n676) );
  or2f U1088 ( .A1(n957), .A2(n956), .Z(n958) );
  or2f U1091 ( .A1(n683), .A2(n921), .Z(n922) );
  inv1f U1092 ( .I(n687), .ZN(n704) );
  or2f U1095 ( .A1(n885), .A2(x1), .Z(n841) );
  and2f U1097 ( .A1(k0), .A2(n788), .Z(n682) );
  and2f U1102 ( .A1(i0), .A2(n788), .Z(n783) );
  or2f U1103 ( .A1(n788), .A2(n787), .Z(n724) );
  or2f U1104 ( .A1(n793), .A2(n792), .Z(n888) );
  and2f U1116 ( .A1(n888), .A2(n681), .Z(n680) );
  inv1f U1129 ( .I(n666), .ZN(n925) );
  and2f U1130 ( .A1(l0), .A2(d2), .Z(n666) );
  and2f U1134 ( .A1(n696), .A2(n697), .Z(n960) );
  or2f U1139 ( .A1(n927), .A2(n926), .Z(n928) );
  or2f U1153 ( .A1(n894), .A2(n893), .Z(n895) );
  and2f U1158 ( .A1(n694), .A2(n891), .Z(n893) );
  or2f U1167 ( .A1(n780), .A2(n804), .Z(n694) );
  inv1f U1168 ( .I(e4), .ZN(n938) );
  or2f U1169 ( .A1(n914), .A2(n913), .Z(n915) );
  or2f U1170 ( .A1(n670), .A2(n915), .Z(n698) );
  and2f U1171 ( .A1(n922), .A2(n702), .Z(n701) );
endmodule

