
module C880_iscas ( h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, 
        s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, 
        a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, 
        d, c, b, a, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, 
        s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1 );
  input h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0,
         p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y,
         x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b,
         a;
  output h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1,
         q1, p1, o1, n1, m1, l1, k1, j1, i1;
  wire   n7, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n107, n108,
         n117, n119, n120, n121, n242, n264, n335, n336, n337, n338, n339,
         n340, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n432,
         n433, n434, n435, n436, n437, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739;

  and2 U4 ( .A1(g1), .A2(c1), .Z(n7) );
  or2 U22 ( .A1(n26), .A2(n27), .Z(y1) );
  inv1 U23 ( .I(n28), .ZN(n27) );
  or2 U24 ( .A1(n29), .A2(n30), .Z(n28) );
  and2 U25 ( .A1(n30), .A2(n29), .Z(n26) );
  and2 U26 ( .A1(n31), .A2(n32), .Z(n29) );
  or2 U27 ( .A1(n33), .A2(u0), .Z(n32) );
  inv1 U28 ( .I(n34), .ZN(n31) );
  and2 U29 ( .A1(n33), .A2(u0), .Z(n34) );
  and2 U30 ( .A1(n35), .A2(n36), .Z(n33) );
  inv1 U31 ( .I(n37), .ZN(n36) );
  and2 U32 ( .A1(n38), .A2(n39), .Z(n37) );
  or2 U33 ( .A1(n39), .A2(n38), .Z(n35) );
  or2 U34 ( .A1(n40), .A2(n41), .Z(n38) );
  and2 U35 ( .A1(n42), .A2(n43), .Z(n41) );
  inv1 U36 ( .I(n44), .ZN(n40) );
  or2 U37 ( .A1(n43), .A2(n42), .Z(n44) );
  or2 U38 ( .A1(n45), .A2(n46), .Z(n42) );
  inv1 U39 ( .I(n47), .ZN(n46) );
  or2 U40 ( .A1(n48), .A2(p0), .Z(n47) );
  and2 U41 ( .A1(p0), .A2(n48), .Z(n45) );
  inv1 U42 ( .I(o0), .ZN(n48) );
  and2 U43 ( .A1(n49), .A2(n50), .Z(n39) );
  inv1 U44 ( .I(n51), .ZN(n50) );
  and2 U45 ( .A1(n52), .A2(n53), .Z(n51) );
  or2 U46 ( .A1(n53), .A2(n52), .Z(n49) );
  or2 U47 ( .A1(n54), .A2(n55), .Z(n52) );
  and2 U48 ( .A1(q0), .A2(n56), .Z(n55) );
  inv1 U49 ( .I(n57), .ZN(n54) );
  or2 U50 ( .A1(n56), .A2(q0), .Z(n57) );
  inv1 U51 ( .I(r0), .ZN(n56) );
  and2 U52 ( .A1(n58), .A2(n59), .Z(n53) );
  or2 U53 ( .A1(n60), .A2(t0), .Z(n59) );
  inv1 U54 ( .I(s0), .ZN(n60) );
  or2 U55 ( .A1(n543), .A2(s0), .Z(n58) );
  or2 U57 ( .A1(n62), .A2(n63), .Z(n30) );
  and2 U58 ( .A1(v0), .A2(n64), .Z(n63) );
  inv1 U59 ( .I(w0), .ZN(n64) );
  and2 U60 ( .A1(w0), .A2(n739), .Z(n62) );
  or2 U62 ( .A1(n65), .A2(n66), .Z(x1) );
  and2 U63 ( .A1(n67), .A2(n68), .Z(n66) );
  inv1 U64 ( .I(n69), .ZN(n65) );
  or2 U65 ( .A1(n68), .A2(n67), .Z(n69) );
  or2 U66 ( .A1(n70), .A2(n71), .Z(n67) );
  inv1 U67 ( .I(n72), .ZN(n71) );
  or2 U68 ( .A1(n73), .A2(d0), .Z(n72) );
  and2 U69 ( .A1(n73), .A2(d0), .Z(n70) );
  and2 U70 ( .A1(n74), .A2(n75), .Z(n73) );
  inv1 U71 ( .I(n76), .ZN(n75) );
  and2 U72 ( .A1(n77), .A2(n78), .Z(n76) );
  or2 U73 ( .A1(n78), .A2(n77), .Z(n74) );
  or2 U74 ( .A1(n79), .A2(n80), .Z(n77) );
  inv1 U75 ( .I(n81), .ZN(n80) );
  or2 U76 ( .A1(n82), .A2(a0), .Z(n81) );
  and2 U77 ( .A1(n82), .A2(a0), .Z(n79) );
  and2 U78 ( .A1(n83), .A2(n84), .Z(n82) );
  or2 U79 ( .A1(n85), .A2(c0), .Z(n84) );
  inv1 U80 ( .I(b0), .ZN(n85) );
  or2 U81 ( .A1(n86), .A2(b0), .Z(n83) );
  inv1 U82 ( .I(c0), .ZN(n86) );
  and2 U83 ( .A1(n87), .A2(n88), .Z(n78) );
  inv1 U84 ( .I(n89), .ZN(n88) );
  and2 U85 ( .A1(n90), .A2(n91), .Z(n89) );
  or2 U86 ( .A1(n91), .A2(n90), .Z(n87) );
  or2 U87 ( .A1(n92), .A2(n93), .Z(n90) );
  inv1 U88 ( .I(n94), .ZN(n93) );
  or2 U89 ( .A1(n43), .A2(x), .Z(n94) );
  and2 U90 ( .A1(x), .A2(n43), .Z(n92) );
  inv1 U91 ( .I(f0), .ZN(n43) );
  and2 U92 ( .A1(n95), .A2(n96), .Z(n91) );
  inv1 U93 ( .I(n97), .ZN(n96) );
  and2 U94 ( .A1(y), .A2(n98), .Z(n97) );
  or2 U95 ( .A1(n98), .A2(y), .Z(n95) );
  inv1 U96 ( .I(z), .ZN(n98) );
  and2 U97 ( .A1(n99), .A2(n100), .Z(n68) );
  or2 U98 ( .A1(n101), .A2(g0), .Z(n100) );
  inv1 U99 ( .I(e0), .ZN(n101) );
  or2 U100 ( .A1(n102), .A2(e0), .Z(n99) );
  inv1 U101 ( .I(g0), .ZN(n102) );
  and2 U102 ( .A1(v), .A2(n103), .Z(w1) );
  and2 U103 ( .A1(n104), .A2(o), .Z(v1) );
  and2 U104 ( .A1(n105), .A2(k), .Z(n104) );
  and2 U105 ( .A1(n105), .A2(f), .Z(u1) );
  inv1 U107 ( .I(k1), .ZN(n107) );
  and2 U108 ( .A1(w), .A2(n103), .Z(r1) );
  or2 U109 ( .A1(t), .A2(u), .Z(n103) );
  inv1 U114 ( .I(g), .ZN(n108) );
  and2 U119 ( .A1(d), .A2(c), .Z(n117) );
  and2 U121 ( .A1(s), .A2(r), .Z(l1) );
  and2 U122 ( .A1(g), .A2(n119), .Z(k1) );
  and2 U123 ( .A1(f), .A2(h), .Z(n119) );
  and2 U124 ( .A1(n120), .A2(g), .Z(j1) );
  and2 U125 ( .A1(q), .A2(f), .Z(n120) );
  and2 U126 ( .A1(n121), .A2(h), .Z(i1) );
  and2 U127 ( .A1(p), .A2(f), .Z(n121) );
  and2 U244 ( .A1(c0), .A2(x0), .Z(n242) );
  and2 U263 ( .A1(b0), .A2(x0), .Z(n264) );
  and2 U359 ( .A1(n), .A2(m), .Z(n336) );
  and2 U360 ( .A1(n105), .A2(n337), .Z(n335) );
  and2 U361 ( .A1(k), .A2(h), .Z(n337) );
  and2 U362 ( .A1(n338), .A2(n339), .Z(n105) );
  and2 U363 ( .A1(c), .A2(l), .Z(n339) );
  and2 U364 ( .A1(b), .A2(n340), .Z(n338) );
  and2 U365 ( .A1(a), .A2(j), .Z(n340) );
  inv1 U371 ( .I(n359), .ZN(n345) );
  inv1 U372 ( .I(n433), .ZN(n346) );
  inv1 U374 ( .I(n347), .ZN(n714) );
  or2 U377 ( .A1(n566), .A2(t0), .Z(n350) );
  or2 U380 ( .A1(n601), .A2(n353), .Z(n352) );
  inv1 U382 ( .I(a1), .ZN(n353) );
  or2 U384 ( .A1(n694), .A2(n693), .Z(n355) );
  or2 U387 ( .A1(n409), .A2(n410), .Z(n358) );
  or2 U388 ( .A1(r0), .A2(n613), .Z(n359) );
  or2 U389 ( .A1(n534), .A2(n360), .Z(n399) );
  or2 U393 ( .A1(n724), .A2(n732), .Z(n362) );
  inv1 U397 ( .I(q0), .ZN(n365) );
  or2 U399 ( .A1(n557), .A2(n369), .Z(n367) );
  or2 U401 ( .A1(n558), .A2(y0), .Z(n368) );
  or2 U402 ( .A1(n586), .A2(n558), .Z(n369) );
  inv1 U405 ( .I(n371), .ZN(n370) );
  or2 U406 ( .A1(n638), .A2(n430), .Z(n372) );
  inv1 U407 ( .I(n372), .ZN(n557) );
  or2 U409 ( .A1(n421), .A2(n375), .Z(n374) );
  inv1 U410 ( .I(n660), .ZN(n375) );
  or2 U411 ( .A1(n650), .A2(n378), .Z(n376) );
  and2 U412 ( .A1(n376), .A2(n377), .Z(e2) );
  or2 U413 ( .A1(n659), .A2(n651), .Z(n377) );
  or2 U414 ( .A1(n649), .A2(n659), .Z(n378) );
  or2 U415 ( .A1(n554), .A2(n382), .Z(n380) );
  and2 U416 ( .A1(n380), .A2(n381), .Z(a2) );
  or2 U417 ( .A1(n556), .A2(n555), .Z(n381) );
  or2 U418 ( .A1(z0), .A2(n556), .Z(n382) );
  or2 U421 ( .A1(n563), .A2(n386), .Z(n384) );
  and2 U422 ( .A1(n384), .A2(n385), .Z(b2) );
  or2 U423 ( .A1(n574), .A2(n564), .Z(n385) );
  or2 U424 ( .A1(n562), .A2(n574), .Z(n386) );
  inv1 U426 ( .I(n387), .ZN(n545) );
  inv1 U428 ( .I(n702), .ZN(n389) );
  inv1 U429 ( .I(n355), .ZN(n390) );
  or2 U430 ( .A1(n373), .A2(n739), .Z(n393) );
  inv1 U436 ( .I(n399), .ZN(n457) );
  inv1 U443 ( .I(f1), .ZN(n405) );
  or2 U446 ( .A1(n409), .A2(n410), .Z(n408) );
  inv1 U448 ( .I(u0), .ZN(n410) );
  or2 U449 ( .A1(n425), .A2(u0), .Z(n411) );
  inv1 U451 ( .I(h), .ZN(n413) );
  and2 U453 ( .A1(n335), .A2(n336), .Z(n415) );
  and2 U462 ( .A1(a), .A2(b), .Z(n422) );
  and2 U465 ( .A1(n703), .A2(y0), .Z(n424) );
  or2 U466 ( .A1(n529), .A2(n528), .Z(n425) );
  or2 U468 ( .A1(n679), .A2(p0), .Z(n427) );
  or2 U469 ( .A1(p0), .A2(n619), .Z(n428) );
  or2 U470 ( .A1(n412), .A2(n739), .Z(n429) );
  and2 U473 ( .A1(n396), .A2(n500), .Z(n432) );
  and2 U475 ( .A1(n605), .A2(r0), .Z(n434) );
  or2 U476 ( .A1(n664), .A2(n665), .Z(n435) );
  or2 U478 ( .A1(n668), .A2(n667), .Z(n436) );
  or2 U479 ( .A1(h1), .A2(n442), .Z(n437) );
  inv1 U481 ( .I(t1), .ZN(n440) );
  inv1 U482 ( .I(n477), .ZN(n441) );
  inv1 U483 ( .I(i), .ZN(n442) );
  or2 U485 ( .A1(n445), .A2(n344), .Z(n444) );
  inv1 U488 ( .I(n486), .ZN(n447) );
  inv1 U490 ( .I(n448), .ZN(n646) );
  inv1 U491 ( .I(d), .ZN(n449) );
  or2 U494 ( .A1(n669), .A2(y0), .Z(n451) );
  or2 U495 ( .A1(n398), .A2(n669), .Z(n452) );
  or2 U496 ( .A1(n407), .A2(n455), .Z(n453) );
  or2 U499 ( .A1(n379), .A2(n419), .Z(n455) );
  and2 U501 ( .A1(n547), .A2(s0), .Z(n458) );
  inv1 U505 ( .I(n460), .ZN(n611) );
  or2 U506 ( .A1(n610), .A2(q0), .Z(n462) );
  inv1 U508 ( .I(n458), .ZN(n637) );
  or2 U509 ( .A1(n467), .A2(n419), .Z(n465) );
  inv1 U511 ( .I(n466), .ZN(n674) );
  inv1 U512 ( .I(y0), .ZN(n467) );
  inv1 U514 ( .I(n445), .ZN(n717) );
  inv1 U515 ( .I(v0), .ZN(n739) );
  inv1 U516 ( .I(a), .ZN(n497) );
  and2 U517 ( .A1(n422), .A2(n117), .Z(m1) );
  inv1 U518 ( .I(e), .ZN(n469) );
  or2 U519 ( .A1(n497), .A2(n469), .Z(n471) );
  inv1 U520 ( .I(n117), .ZN(n470) );
  or2 U521 ( .A1(n471), .A2(n470), .Z(n476) );
  or2 U522 ( .A1(n476), .A2(k1), .Z(n1) );
  inv1 U523 ( .I(p), .ZN(n472) );
  inv1 U524 ( .I(q), .ZN(n473) );
  or2 U525 ( .A1(n472), .A2(n473), .Z(n479) );
  inv1 U526 ( .I(k), .ZN(n491) );
  or2 U527 ( .A1(n479), .A2(n491), .Z(o1) );
  or2 U528 ( .A1(n473), .A2(n491), .Z(n474) );
  or2 U529 ( .A1(n474), .A2(n108), .Z(p1) );
  inv1 U530 ( .I(h), .ZN(n487) );
  or2 U531 ( .A1(n491), .A2(n487), .Z(n475) );
  or2 U532 ( .A1(n475), .A2(n108), .Z(q1) );
  or2 U533 ( .A1(n476), .A2(n107), .Z(s1) );
  and2 U535 ( .A1(y0), .A2(n405), .Z(n503) );
  or2 U536 ( .A1(n437), .A2(n441), .Z(n481) );
  inv1 U537 ( .I(f), .ZN(n478) );
  inv1 U540 ( .I(j), .ZN(n482) );
  and2 U545 ( .A1(i), .A2(d), .Z(n484) );
  or2 U547 ( .A1(n413), .A2(d), .Z(n489) );
  inv1 U550 ( .I(n0), .ZN(n490) );
  and2 U557 ( .A1(i), .A2(e), .Z(n495) );
  and2 U558 ( .A1(n495), .A2(d), .Z(n496) );
  or2 U562 ( .A1(n373), .A2(n739), .Z(n500) );
  or2 U565 ( .A1(n627), .A2(n501), .Z(n504) );
  or2 U567 ( .A1(n503), .A2(n502), .Z(n508) );
  and2 U568 ( .A1(y0), .A2(f1), .Z(n506) );
  inv1 U569 ( .I(n504), .ZN(n505) );
  or2 U570 ( .A1(n506), .A2(n505), .Z(n507) );
  and2 U571 ( .A1(n508), .A2(n507), .Z(n510) );
  and2 U572 ( .A1(x0), .A2(d0), .Z(n509) );
  or2 U573 ( .A1(n510), .A2(n509), .Z(n511) );
  or2 U574 ( .A1(n511), .A2(n7), .Z(n518) );
  and2 U575 ( .A1(b1), .A2(n392), .Z(n516) );
  and2 U576 ( .A1(v0), .A2(n415), .Z(n514) );
  and2 U577 ( .A1(a1), .A2(n627), .Z(n513) );
  or2 U578 ( .A1(n514), .A2(n513), .Z(n515) );
  or2 U579 ( .A1(n516), .A2(n515), .Z(n517) );
  or2 U580 ( .A1(n518), .A2(n517), .Z(z1) );
  and2 U581 ( .A1(i0), .A2(n530), .Z(n520) );
  and2 U584 ( .A1(a1), .A2(n458), .Z(n526) );
  and2 U585 ( .A1(b1), .A2(n547), .Z(n524) );
  and2 U586 ( .A1(s0), .A2(n415), .Z(n522) );
  and2 U587 ( .A1(a0), .A2(x0), .Z(n521) );
  or2 U588 ( .A1(n522), .A2(n521), .Z(n523) );
  or2 U589 ( .A1(n524), .A2(n523), .Z(n525) );
  or2 U590 ( .A1(n526), .A2(n525), .Z(n556) );
  inv1 U596 ( .I(n687), .ZN(n638) );
  or2 U607 ( .A1(n540), .A2(n541), .Z(n542) );
  inv1 U609 ( .I(n566), .ZN(n544) );
  inv1 U610 ( .I(t0), .ZN(n543) );
  or2 U611 ( .A1(n544), .A2(n543), .Z(n695) );
  inv1 U613 ( .I(n358), .ZN(n586) );
  and2 U615 ( .A1(y0), .A2(n550), .Z(n549) );
  or2 U616 ( .A1(n458), .A2(n366), .Z(n552) );
  inv1 U617 ( .I(n552), .ZN(n548) );
  or2 U618 ( .A1(n549), .A2(n548), .Z(n555) );
  inv1 U619 ( .I(n550), .ZN(n551) );
  and2 U620 ( .A1(y0), .A2(n551), .Z(n553) );
  or2 U621 ( .A1(n553), .A2(n552), .Z(n554) );
  or2 U622 ( .A1(n557), .A2(n586), .Z(n559) );
  or2 U623 ( .A1(n567), .A2(n691), .Z(n561) );
  inv1 U624 ( .I(n561), .ZN(n558) );
  inv1 U625 ( .I(n559), .ZN(n560) );
  or2 U627 ( .A1(n561), .A2(z0), .Z(n562) );
  and2 U628 ( .A1(d1), .A2(c1), .Z(n565) );
  or2 U629 ( .A1(n565), .A2(n264), .Z(n573) );
  and2 U630 ( .A1(t0), .A2(n415), .Z(n571) );
  and2 U631 ( .A1(b1), .A2(n566), .Z(n569) );
  or2 U633 ( .A1(n569), .A2(n568), .Z(n570) );
  or2 U634 ( .A1(n571), .A2(n570), .Z(n572) );
  or2 U635 ( .A1(n573), .A2(n572), .Z(n574) );
  and2 U636 ( .A1(y0), .A2(n430), .Z(n576) );
  or2 U638 ( .A1(n577), .A2(z0), .Z(n575) );
  or2 U639 ( .A1(n576), .A2(n575), .Z(n581) );
  and2 U640 ( .A1(y0), .A2(n400), .Z(n579) );
  inv1 U641 ( .I(n577), .ZN(n578) );
  or2 U642 ( .A1(n579), .A2(n578), .Z(n580) );
  and2 U643 ( .A1(n581), .A2(n580), .Z(n583) );
  and2 U644 ( .A1(e1), .A2(c1), .Z(n582) );
  or2 U646 ( .A1(n584), .A2(n242), .Z(n592) );
  and2 U647 ( .A1(u0), .A2(n415), .Z(n590) );
  and2 U648 ( .A1(b1), .A2(n425), .Z(n588) );
  and2 U649 ( .A1(a1), .A2(n586), .Z(n587) );
  or2 U650 ( .A1(n588), .A2(n587), .Z(n589) );
  or2 U651 ( .A1(n590), .A2(n589), .Z(n591) );
  or2 U652 ( .A1(n592), .A2(n591), .Z(c2) );
  and2 U653 ( .A1(h0), .A2(b), .Z(n594) );
  and2 U658 ( .A1(i0), .A2(n617), .Z(n598) );
  or2 U659 ( .A1(n598), .A2(n417), .Z(n599) );
  and2 U662 ( .A1(l0), .A2(h0), .Z(n604) );
  and2 U666 ( .A1(h0), .A2(d), .Z(n606) );
  and2 U669 ( .A1(k0), .A2(n617), .Z(n607) );
  or2 U670 ( .A1(n608), .A2(n607), .Z(n609) );
  or2 U672 ( .A1(n407), .A2(n379), .Z(n623) );
  or2 U673 ( .A1(n433), .A2(n613), .Z(n654) );
  and2 U675 ( .A1(h0), .A2(i), .Z(n616) );
  or2 U677 ( .A1(n615), .A2(n616), .Z(n620) );
  and2 U678 ( .A1(j0), .A2(n617), .Z(n618) );
  or2 U679 ( .A1(n618), .A2(n417), .Z(n619) );
  or2 U681 ( .A1(n428), .A2(n620), .Z(n684) );
  and2 U684 ( .A1(n696), .A2(n684), .Z(n624) );
  and2 U690 ( .A1(n632), .A2(n357), .Z(n633) );
  or2 U693 ( .A1(n663), .A2(o0), .Z(n660) );
  and2 U694 ( .A1(n670), .A2(n660), .Z(n636) );
  or2 U695 ( .A1(n421), .A2(n636), .Z(d2) );
  and2 U696 ( .A1(y0), .A2(n637), .Z(n641) );
  or2 U697 ( .A1(n457), .A2(n638), .Z(n639) );
  or2 U698 ( .A1(n366), .A2(n639), .Z(n640) );
  or2 U703 ( .A1(n648), .A2(z0), .Z(n643) );
  or2 U704 ( .A1(n644), .A2(n643), .Z(n651) );
  and2 U706 ( .A1(y0), .A2(n647), .Z(n650) );
  inv1 U707 ( .I(n648), .ZN(n649) );
  and2 U708 ( .A1(z), .A2(x0), .Z(n653) );
  and2 U709 ( .A1(r0), .A2(n415), .Z(n652) );
  or2 U710 ( .A1(n653), .A2(n652), .Z(n658) );
  and2 U711 ( .A1(b1), .A2(n654), .Z(n656) );
  and2 U712 ( .A1(a1), .A2(n434), .Z(n655) );
  or2 U713 ( .A1(n656), .A2(n655), .Z(n657) );
  or2 U714 ( .A1(n658), .A2(n657), .Z(n659) );
  inv1 U715 ( .I(n374), .ZN(n668) );
  and2 U716 ( .A1(x0), .A2(h1), .Z(n662) );
  and2 U717 ( .A1(o0), .A2(n415), .Z(n661) );
  or2 U718 ( .A1(n662), .A2(n661), .Z(n667) );
  and2 U719 ( .A1(b1), .A2(n663), .Z(n665) );
  or2 U721 ( .A1(n667), .A2(n666), .Z(n671) );
  or2 U722 ( .A1(n374), .A2(n671), .Z(n672) );
  or2 U723 ( .A1(n672), .A2(z0), .Z(n673) );
  or2 U724 ( .A1(n674), .A2(n673), .Z(n675) );
  and2 U725 ( .A1(n676), .A2(n675), .Z(f2) );
  and2 U726 ( .A1(x), .A2(x0), .Z(n678) );
  and2 U727 ( .A1(p0), .A2(n415), .Z(n677) );
  or2 U728 ( .A1(n678), .A2(n677), .Z(n683) );
  and2 U729 ( .A1(b1), .A2(n679), .Z(n681) );
  and2 U730 ( .A1(a1), .A2(n419), .Z(n680) );
  or2 U731 ( .A1(n681), .A2(n680), .Z(n682) );
  inv1 U733 ( .I(n427), .ZN(n685) );
  or2 U734 ( .A1(n685), .A2(n419), .Z(n706) );
  or2 U735 ( .A1(z0), .A2(n706), .Z(n686) );
  or2 U736 ( .A1(n708), .A2(n686), .Z(n705) );
  inv1 U741 ( .I(n350), .ZN(n691) );
  or2 U742 ( .A1(n691), .A2(n366), .Z(n692) );
  or2 U744 ( .A1(n694), .A2(n693), .Z(n703) );
  or2 U749 ( .A1(n611), .A2(n406), .Z(n700) );
  inv1 U751 ( .I(n706), .ZN(n707) );
  or2 U752 ( .A1(n708), .A2(n707), .Z(n709) );
  or2 U753 ( .A1(n423), .A2(n709), .Z(n710) );
  and2 U754 ( .A1(n710), .A2(n711), .Z(g2) );
  inv1 U758 ( .I(n729), .ZN(n716) );
  and2 U759 ( .A1(y0), .A2(n716), .Z(n718) );
  or2 U762 ( .A1(n379), .A2(n697), .Z(n732) );
  and2 U763 ( .A1(y), .A2(x0), .Z(n720) );
  and2 U764 ( .A1(q0), .A2(n415), .Z(n719) );
  or2 U765 ( .A1(n720), .A2(n719), .Z(n724) );
  and2 U766 ( .A1(b1), .A2(n416), .Z(n722) );
  and2 U767 ( .A1(a1), .A2(n379), .Z(n721) );
  or2 U768 ( .A1(n722), .A2(n721), .Z(n723) );
  or2 U769 ( .A1(n724), .A2(n723), .Z(n733) );
  or2 U770 ( .A1(n723), .A2(n362), .Z(n725) );
  or2 U771 ( .A1(n725), .A2(z0), .Z(n726) );
  or2 U772 ( .A1(n727), .A2(n726), .Z(n738) );
  inv1 U773 ( .I(n728), .ZN(n730) );
  inv1 U776 ( .I(n732), .ZN(n734) );
  or2 U777 ( .A1(n734), .A2(n733), .Z(n735) );
  or2 U778 ( .A1(n736), .A2(n735), .Z(n737) );
  and2 U779 ( .A1(n738), .A2(n737), .Z(h2) );
  inv1f U366 ( .I(n696), .ZN(n697) );
  inv1f U367 ( .I(n344), .ZN(n391) );
  or2f U368 ( .A1(n461), .A2(n633), .Z(n670) );
  and2f U369 ( .A1(n453), .A2(n454), .Z(n461) );
  or2 U370 ( .A1(n491), .A2(n490), .Z(n595) );
  and2 U373 ( .A1(n447), .A2(n485), .Z(n446) );
  and2 U375 ( .A1(m0), .A2(n617), .Z(n603) );
  inv1 U376 ( .I(n536), .ZN(n531) );
  or2 U378 ( .A1(n504), .A2(z0), .Z(n502) );
  inv1 U379 ( .I(n429), .ZN(n627) );
  inv1 U381 ( .I(n392), .ZN(n412) );
  or2f U383 ( .A1(n499), .A2(n383), .Z(n392) );
  and2f U385 ( .A1(n361), .A2(n391), .Z(n713) );
  or2f U386 ( .A1(n379), .A2(n391), .Z(n621) );
  or2f U390 ( .A1(n698), .A2(n697), .Z(n699) );
  or2f U391 ( .A1(n344), .A2(n697), .Z(n406) );
  or2f U392 ( .A1(n697), .A2(n688), .Z(n689) );
  and2f U394 ( .A1(n424), .A2(n702), .Z(n704) );
  and2f U395 ( .A1(n679), .A2(p0), .Z(n419) );
  or2f U396 ( .A1(n620), .A2(n619), .Z(n679) );
  inv1 U398 ( .I(n512), .ZN(n373) );
  inv1 U400 ( .I(n585), .ZN(n409) );
  or2 U403 ( .A1(n434), .A2(n344), .Z(n648) );
  or2 U404 ( .A1(n699), .A2(n344), .Z(n701) );
  or2 U408 ( .A1(n449), .A2(h), .Z(n488) );
  and2 U419 ( .A1(k), .A2(p), .Z(n483) );
  and2 U420 ( .A1(n538), .A2(a0), .Z(n414) );
  inv1 U425 ( .I(n393), .ZN(n401) );
  or2 U427 ( .A1(n688), .A2(n586), .Z(n577) );
  inv1 U431 ( .I(n597), .ZN(n418) );
  and2 U432 ( .A1(n614), .A2(z), .Z(n608) );
  and2 U433 ( .A1(n614), .A2(d0), .Z(n394) );
  or2 U434 ( .A1(n604), .A2(n603), .Z(n613) );
  or2 U435 ( .A1(n414), .A2(n417), .Z(n433) );
  and2 U437 ( .A1(n614), .A2(b0), .Z(n519) );
  and2 U438 ( .A1(y), .A2(n614), .Z(n615) );
  and2 U439 ( .A1(n628), .A2(n629), .Z(n630) );
  and2 U440 ( .A1(n623), .A2(n622), .Z(n634) );
  or2 U441 ( .A1(n690), .A2(n689), .Z(n694) );
  and2 U442 ( .A1(n629), .A2(n628), .Z(n348) );
  and2 U444 ( .A1(n641), .A2(n645), .Z(n642) );
  or2 U445 ( .A1(n717), .A2(n448), .Z(n647) );
  and2 U447 ( .A1(n367), .A2(n368), .Z(n564) );
  or2 U450 ( .A1(n704), .A2(n705), .Z(n711) );
  inv1 U452 ( .I(n400), .ZN(n430) );
  or2f U454 ( .A1(n401), .A2(n402), .Z(n400) );
  inv1 U455 ( .I(n396), .ZN(n402) );
  inv1 U456 ( .I(n361), .ZN(n366) );
  and2 U457 ( .A1(n695), .A2(n387), .Z(n347) );
  inv1 U458 ( .I(n364), .ZN(n379) );
  inv1f U459 ( .I(n352), .ZN(n664) );
  and2f U460 ( .A1(n718), .A2(n444), .Z(n727) );
  and2 U461 ( .A1(n426), .A2(n361), .Z(n448) );
  and2f U463 ( .A1(y0), .A2(n560), .Z(n563) );
  or2f U464 ( .A1(n394), .A2(n395), .Z(n687) );
  or2f U467 ( .A1(n397), .A2(n634), .Z(n635) );
  or2f U471 ( .A1(n635), .A2(n465), .Z(n466) );
  or2f U472 ( .A1(n493), .A2(n440), .Z(n494) );
  and2f U474 ( .A1(n739), .A2(n373), .Z(n501) );
  or2f U477 ( .A1(n499), .A2(n354), .Z(n512) );
  and2f U480 ( .A1(n500), .A2(n396), .Z(n349) );
  and2f U484 ( .A1(e), .A2(a), .Z(n477) );
  or2f U486 ( .A1(n608), .A2(n363), .Z(n416) );
  or2f U487 ( .A1(n610), .A2(n607), .Z(n363) );
  or2f U489 ( .A1(n683), .A2(n682), .Z(n708) );
  or2f U492 ( .A1(n665), .A2(n664), .Z(n666) );
  inv1f U493 ( .I(n421), .ZN(n601) );
  and2f U497 ( .A1(h), .A2(n483), .Z(n486) );
  or2f U498 ( .A1(n714), .A2(n546), .Z(n550) );
  and2f U500 ( .A1(n400), .A2(n629), .Z(n546) );
  and2f U502 ( .A1(n422), .A2(n484), .Z(n485) );
  inv1f U503 ( .I(n536), .ZN(n537) );
  or2f U504 ( .A1(t0), .A2(n537), .Z(n351) );
  and2f U507 ( .A1(n645), .A2(n637), .Z(n445) );
  or2f U510 ( .A1(n606), .A2(n417), .Z(n610) );
  and2f U513 ( .A1(n391), .A2(n624), .Z(n625) );
  or2f U534 ( .A1(n462), .A2(n609), .Z(n696) );
  or2f U538 ( .A1(n529), .A2(n528), .Z(n585) );
  and2f U539 ( .A1(n642), .A2(n646), .Z(n644) );
  or2f U541 ( .A1(n567), .A2(n545), .Z(n426) );
  or2f U542 ( .A1(n366), .A2(n695), .Z(n698) );
  and2f U543 ( .A1(a1), .A2(n567), .Z(n568) );
  inv1f U544 ( .I(n695), .ZN(n567) );
  or2f U546 ( .A1(n351), .A2(n532), .Z(n360) );
  or2f U548 ( .A1(n532), .A2(n537), .Z(n533) );
  and2f U549 ( .A1(k0), .A2(n530), .Z(n527) );
  and2f U551 ( .A1(j0), .A2(n530), .Z(n532) );
  or2f U552 ( .A1(n531), .A2(n420), .Z(n354) );
  or2f U553 ( .A1(n420), .A2(n531), .Z(n383) );
  or2f U554 ( .A1(n531), .A2(n420), .Z(n541) );
  and2f U555 ( .A1(n450), .A2(n451), .Z(n676) );
  or2f U556 ( .A1(n452), .A2(n461), .Z(n450) );
  and2f U559 ( .A1(n538), .A2(e0), .Z(n539) );
  and2f U560 ( .A1(n343), .A2(i), .Z(t1) );
  and2f U561 ( .A1(e), .A2(a), .Z(n343) );
  and2f U563 ( .A1(n614), .A2(d0), .Z(n529) );
  and2f U564 ( .A1(n614), .A2(e0), .Z(n499) );
  and2f U566 ( .A1(x), .A2(n614), .Z(n593) );
  and2f U582 ( .A1(n388), .A2(y0), .Z(n423) );
  or2f U583 ( .A1(n389), .A2(n390), .Z(n388) );
  and2f U591 ( .A1(n496), .A2(n595), .Z(n498) );
  or2f U592 ( .A1(n519), .A2(n443), .Z(n547) );
  or2f U593 ( .A1(n531), .A2(n520), .Z(n443) );
  or2f U594 ( .A1(n547), .A2(s0), .Z(n361) );
  or2f U595 ( .A1(n612), .A2(n613), .Z(n605) );
  or2f U597 ( .A1(n414), .A2(n417), .Z(n612) );
  and2f U598 ( .A1(n621), .A2(n427), .Z(n622) );
  and2f U599 ( .A1(n460), .A2(n696), .Z(n407) );
  or2f U600 ( .A1(n531), .A2(n527), .Z(n528) );
  or2f U601 ( .A1(n527), .A2(n370), .Z(n395) );
  or2f U602 ( .A1(n688), .A2(n457), .Z(n535) );
  inv1f U603 ( .I(n411), .ZN(n688) );
  or2f U604 ( .A1(n539), .A2(v0), .Z(n540) );
  or2f U605 ( .A1(n583), .A2(n582), .Z(n584) );
  or2f U606 ( .A1(n492), .A2(n595), .Z(n493) );
  and2f U608 ( .A1(n731), .A2(y0), .Z(n736) );
  or2f U612 ( .A1(n730), .A2(n729), .Z(n731) );
  or2f U614 ( .A1(n715), .A2(n434), .Z(n729) );
  and2f U626 ( .A1(n426), .A2(n713), .Z(n715) );
  or2f U632 ( .A1(n534), .A2(n533), .Z(n566) );
  and2f U637 ( .A1(n538), .A2(c0), .Z(n534) );
  and2f U645 ( .A1(n645), .A2(n637), .Z(n468) );
  and2f U654 ( .A1(n536), .A2(n410), .Z(n371) );
  or2f U655 ( .A1(n432), .A2(n640), .Z(n645) );
  or2f U656 ( .A1(n597), .A2(n482), .Z(n536) );
  and2f U657 ( .A1(n349), .A2(n358), .Z(n690) );
  or2f U660 ( .A1(n404), .A2(n405), .Z(n396) );
  inv1f U661 ( .I(n542), .ZN(n404) );
  or2f U663 ( .A1(n498), .A2(n497), .Z(n530) );
  and2f U664 ( .A1(n530), .A2(m0), .Z(n420) );
  or2f U665 ( .A1(n435), .A2(n436), .Z(n669) );
  or2f U667 ( .A1(n600), .A2(n599), .Z(n663) );
  or2f U668 ( .A1(n594), .A2(n593), .Z(n600) );
  and2f U671 ( .A1(n663), .A2(o0), .Z(n421) );
  or2f U674 ( .A1(n602), .A2(n446), .Z(n614) );
  or2f U676 ( .A1(n456), .A2(n464), .Z(n460) );
  and2f U680 ( .A1(n547), .A2(s0), .Z(n464) );
  and2f U682 ( .A1(n605), .A2(r0), .Z(n456) );
  and2f U683 ( .A1(n459), .A2(n701), .Z(n702) );
  and2f U685 ( .A1(n700), .A2(n364), .Z(n459) );
  and2f U686 ( .A1(n596), .A2(n595), .Z(n617) );
  and2f U687 ( .A1(t1), .A2(j), .Z(n596) );
  and2f U688 ( .A1(n357), .A2(n632), .Z(n398) );
  or2f U689 ( .A1(n348), .A2(n714), .Z(n357) );
  or2f U691 ( .A1(n408), .A2(n691), .Z(n387) );
  or2f U692 ( .A1(n481), .A2(n480), .Z(n597) );
  or2f U699 ( .A1(n479), .A2(n478), .Z(n480) );
  or2f U700 ( .A1(n419), .A2(n622), .Z(n454) );
  or2f U701 ( .A1(n463), .A2(n365), .Z(n364) );
  inv1f U702 ( .I(n416), .ZN(n463) );
  and2f U705 ( .A1(n418), .A2(d), .Z(n417) );
  or2f U720 ( .A1(n692), .A2(n344), .Z(n693) );
  or2f U732 ( .A1(n468), .A2(n344), .Z(n728) );
  and2f U737 ( .A1(n345), .A2(n346), .Z(n344) );
  inv1f U738 ( .I(n535), .ZN(n629) );
  or2f U739 ( .A1(n627), .A2(n402), .Z(n628) );
  and2f U740 ( .A1(n631), .A2(n632), .Z(n397) );
  and2f U743 ( .A1(n625), .A2(n361), .Z(n632) );
  or2f U745 ( .A1(n630), .A2(n714), .Z(n631) );
  and2f U746 ( .A1(n489), .A2(n488), .Z(n492) );
  or2f U747 ( .A1(n602), .A2(n446), .Z(n538) );
  inv1f U748 ( .I(n494), .ZN(n602) );
endmodule

