
module rot ( e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, 
        o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, y2, x2, 
        w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, g2, f2, 
        e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, 
        m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, 
        u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, 
        c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, 
        f, e, d, c, b, a, h8, g8, f8, e8, d8, c8, b8, a8, z7, y7, x7, w7, v7, 
        u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, 
        c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, 
        k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, 
        s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, 
        a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, 
        i4, h4, g4, f4 );
  input e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3,
         m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, y2, x2, w2,
         v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, g2, f2,
         e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1,
         n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0,
         w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0,
         f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l,
         k, j, i, h, g, f, e, d, c, b, a;
  output h8, g8, f8, e8, d8, c8, b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7,
         q7, p7, o7, n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7,
         z6, y6, x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6,
         i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, s5,
         r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5,
         a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4,
         j4, i4, h4, g4, f4;
  wire   n940, n941, n942, n943, n944, n945, n124, n126, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n158,
         n159, n160, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n183, n184, n205, n206, n207,
         n208, n209, n211, n212, n222, n224, n226, n235, n239, n240, n241,
         n242, n243, n244, n246, n249, n250, n251, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n288, n289, n290, n291, n292, n303, n304,
         n317, n318, n319, n320, n321, n322, n346, n347, n349, n350, n351,
         n352, n353, n354, n355, n356, n360, n362, n363, n364, n365, n366,
         n367, n375, n376, n377, n378, n379, n380, n387, n389, n390, n391,
         n392, n393, n394, n395, n396, n399, n400, n402, n403, n404, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n422, n423, n424, n425, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n458, n459, n467, n477, n478, n479, n480, n481, n482, n484,
         n486, n487, n488, n489, n490, n491, n495, n496, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n520, n521, n522, n526,
         n527, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n611, n613, n614,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n647, n648, n649, n650, n651, n653, n655, n656, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n717, n718, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n785, n786, n787, n788, n790, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n841, n842, n843, n844, n845, n846, n847, n848, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n922, n923, n924, n925, n927, n928, n929, n930, n931, n932,
         n934, n935, n936, n937, n938, n939, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003;

  or2f U241 ( .A1(n390), .A2(n363), .Z(n389) );
  or2f U242 ( .A1(n391), .A2(n392), .Z(n363) );
  and2f U243 ( .A1(n393), .A2(n394), .Z(n392) );
  or2f U281 ( .A1(n425), .A2(n428), .Z(n427) );
  and2f U282 ( .A1(n393), .A2(n429), .Z(n428) );
  or2f U283 ( .A1(n979), .A2(n395), .Z(n429) );
  or2f U554 ( .A1(n924), .A2(g2), .Z(n379) );
  or2f U556 ( .A1(n617), .A2(n320), .Z(n264) );
  and2f U612 ( .A1(x1), .A2(m2), .Z(n173) );
  and2f U619 ( .A1(n303), .A2(n304), .Z(n651) );
  and2f U626 ( .A1(n173), .A2(y1), .Z(n655) );
  buf0 U629 ( .I(n935), .Z(h4) );
  buf0 U630 ( .I(n934), .Z(i4) );
  buf0 U631 ( .I(n931), .Z(j4) );
  buf0 U632 ( .I(s3), .Z(k4) );
  buf0 U633 ( .I(n945), .Z(l4) );
  buf0 U634 ( .I(t3), .Z(m4) );
  buf0 U635 ( .I(m2), .Z(a5) );
  buf0 U636 ( .I(l2), .Z(k5) );
  buf0 U637 ( .I(n944), .Z(d6) );
  buf0 U638 ( .I(n943), .Z(k6) );
  buf0 U639 ( .I(n941), .Z(v6) );
  buf0 U640 ( .I(y0), .Z(w6) );
  buf0 U641 ( .I(n942), .Z(x6) );
  buf0 U642 ( .I(w0), .Z(y6) );
  buf0 U643 ( .I(n941), .Z(z6) );
  buf0 U644 ( .I(y0), .Z(a7) );
  buf0 U645 ( .I(z0), .Z(b7) );
  buf0 U646 ( .I(n940), .Z(i7) );
  buf0 U647 ( .I(w), .Z(s7) );
  buf0 U648 ( .I(z), .Z(t7) );
  buf0 U649 ( .I(a0), .Z(u7) );
  buf0 U650 ( .I(b0), .Z(v7) );
  buf0 U651 ( .I(c0), .Z(w7) );
  buf0 U652 ( .I(n932), .Z(d8) );
  buf0 U653 ( .I(n942), .Z(e8) );
  buf0 U654 ( .I(w0), .Z(f8) );
  buf0 U655 ( .I(x0), .Z(g8) );
  or2 U659 ( .A1(n684), .A2(n881), .Z(n882) );
  and2 U660 ( .A1(n886), .A2(n1000), .Z(n888) );
  and2f U662 ( .A1(n768), .A2(n687), .Z(n685) );
  or2f U663 ( .A1(n685), .A2(n686), .Z(n692) );
  and2f U664 ( .A1(n998), .A2(n771), .Z(n686) );
  or2f U667 ( .A1(n688), .A2(n689), .Z(n750) );
  and2f U668 ( .A1(y3), .A2(n748), .Z(n689) );
  inv1 U671 ( .I(n691), .ZN(n932) );
  and2 U673 ( .A1(a4), .A2(n955), .Z(n910) );
  and2 U675 ( .A1(n887), .A2(n684), .Z(n7) );
  and2 U676 ( .A1(n887), .A2(n1000), .Z(n884) );
  inv1 U677 ( .I(n887), .ZN(n895) );
  or2 U678 ( .A1(n932), .A2(m1), .Z(n879) );
  or2 U679 ( .A1(n932), .A2(n916), .Z(n917) );
  and2 U680 ( .A1(i0), .A2(n868), .Z(n792) );
  or2 U681 ( .A1(n932), .A2(z3), .Z(n850) );
  or2 U682 ( .A1(n932), .A2(v2), .Z(n935) );
  or2 U683 ( .A1(n868), .A2(n354), .Z(n741) );
  or2f U688 ( .A1(n379), .A2(n264), .Z(n873) );
  and2f U689 ( .A1(n782), .A2(n873), .Z(n693) );
  or2f U691 ( .A1(n693), .A2(n803), .Z(n694) );
  or2f U692 ( .A1(n695), .A2(n694), .Z(n467) );
  or2f U714 ( .A1(n701), .A2(n427), .Z(n303) );
  and2f U720 ( .A1(u), .A2(s0), .Z(n703) );
  or2f U734 ( .A1(n911), .A2(n707), .Z(n710) );
  or2f U736 ( .A1(n708), .A2(d0), .Z(n709) );
  or2f U738 ( .A1(n711), .A2(n712), .Z(n715) );
  or2f U741 ( .A1(n715), .A2(n714), .Z(n728) );
  and2f U745 ( .A1(n729), .A2(x2), .Z(n721) );
  inv1f U748 ( .I(k), .ZN(n717) );
  and2f U749 ( .A1(d0), .A2(n717), .Z(n718) );
  or2f U750 ( .A1(n718), .A2(n963), .Z(n720) );
  and2f U751 ( .A1(n720), .A2(n721), .Z(n724) );
  or2f U754 ( .A1(n724), .A2(n723), .Z(n725) );
  and2f U755 ( .A1(n725), .A2(n726), .Z(n727) );
  or2f U756 ( .A1(n727), .A2(n728), .Z(n732) );
  or2f U783 ( .A1(n746), .A2(n932), .Z(n934) );
  or2f U789 ( .A1(n750), .A2(n893), .Z(n890) );
  inv1f U790 ( .I(n890), .ZN(n756) );
  or2f U796 ( .A1(n756), .A2(n755), .Z(n898) );
  and2f U801 ( .A1(n983), .A2(n761), .Z(n813) );
  and2f U804 ( .A1(n983), .A2(n763), .Z(n811) );
  or2f U805 ( .A1(n813), .A2(n811), .Z(n794) );
  and2f U806 ( .A1(n794), .A2(n999), .Z(n765) );
  or2f U807 ( .A1(n765), .A2(n898), .Z(n766) );
  and2f U808 ( .A1(n766), .A2(n955), .Z(n768) );
  and2f U821 ( .A1(n1003), .A2(n998), .Z(n781) );
  inv1f U836 ( .I(n935), .ZN(n795) );
  and2f U837 ( .A1(n934), .A2(n795), .Z(n798) );
  and2f U838 ( .A1(n796), .A2(n935), .Z(n797) );
  or2f U839 ( .A1(n798), .A2(n797), .Z(n814) );
  or2f U840 ( .A1(n799), .A2(n814), .Z(n800) );
  or2f U841 ( .A1(n801), .A2(n800), .Z(n802) );
  and2f U842 ( .A1(n957), .A2(n802), .Z(n810) );
  and2f U851 ( .A1(n988), .A2(n808), .Z(n809) );
  or2f U852 ( .A1(n810), .A2(n809), .Z(t4) );
  and2f U856 ( .A1(n957), .A2(n816), .Z(n819) );
  and2f U858 ( .A1(n988), .A2(n817), .Z(n818) );
  or2f U859 ( .A1(n819), .A2(n818), .Z(u4) );
  and2f U864 ( .A1(d2), .A2(n989), .Z(n833) );
  and2f U869 ( .A1(n988), .A2(n831), .Z(n832) );
  or2f U870 ( .A1(n833), .A2(n832), .Z(w4) );
  and2f U871 ( .A1(e2), .A2(n957), .Z(n842) );
  and2f U877 ( .A1(n988), .A2(n839), .Z(n841) );
  or2f U878 ( .A1(n842), .A2(n841), .Z(x4) );
  and2f U880 ( .A1(n902), .A2(n844), .Z(n846) );
  inv1f U887 ( .I(n863), .ZN(n853) );
  and2f U894 ( .A1(n861), .A2(n860), .Z(q5) );
  and2f U898 ( .A1(n867), .A2(n866), .Z(r5) );
  or2f U901 ( .A1(n870), .A2(n869), .Z(n871) );
  and2f U902 ( .A1(l0), .A2(n871), .Z(n872) );
  or2f U903 ( .A1(n872), .A2(z1), .Z(n875) );
  and2f U911 ( .A1(u2), .A2(n989), .Z(n883) );
  or2f U914 ( .A1(n883), .A2(n882), .Z(l7) );
  and2f U920 ( .A1(n684), .A2(n892), .Z(n897) );
  or2f U921 ( .A1(n893), .A2(n998), .Z(n894) );
  and2f U922 ( .A1(n895), .A2(n894), .Z(n896) );
  or2f U923 ( .A1(n897), .A2(n896), .Z(n908) );
  and2f U925 ( .A1(n1000), .A2(n899), .Z(n901) );
  and2f U929 ( .A1(n906), .A2(n905), .Z(n907) );
  or2f U930 ( .A1(n908), .A2(n907), .Z(n909) );
  and2f U931 ( .A1(n910), .A2(n909), .Z(p7) );
  inv1f U620 ( .I(h0), .ZN(n971) );
  inv1 U621 ( .I(j), .ZN(n707) );
  or2 U622 ( .A1(n998), .A2(n891), .Z(n892) );
  or2 U623 ( .A1(n875), .A2(n874), .Z(u5) );
  or2 U624 ( .A1(n985), .A2(n946), .Z(n776) );
  or2 U625 ( .A1(n986), .A2(n735), .Z(n946) );
  and2f U627 ( .A1(n710), .A2(n709), .Z(n711) );
  inv1f U628 ( .I(n984), .ZN(n1001) );
  and2 U656 ( .A1(n613), .A2(n614), .Z(n611) );
  or2 U657 ( .A1(r1), .A2(n288), .Z(n614) );
  and2 U658 ( .A1(n759), .A2(n758), .Z(n760) );
  and2 U661 ( .A1(u3), .A2(n722), .Z(n723) );
  inv1 U665 ( .I(h), .ZN(n722) );
  and2 U666 ( .A1(u3), .A2(n713), .Z(n714) );
  inv1 U669 ( .I(i), .ZN(n713) );
  or2 U670 ( .A1(n778), .A2(n777), .Z(n820) );
  and2 U672 ( .A1(n959), .A2(n960), .Z(n864) );
  or2 U674 ( .A1(n846), .A2(n961), .Z(n959) );
  inv1 U684 ( .I(g3), .ZN(n978) );
  inv1 U685 ( .I(l), .ZN(n708) );
  inv1 U686 ( .I(g), .ZN(n712) );
  and2 U687 ( .A1(m3), .A2(n400), .Z(n762) );
  and2 U690 ( .A1(x2), .A2(n728), .Z(n981) );
  inv1 U693 ( .I(n934), .ZN(n796) );
  and2 U694 ( .A1(n774), .A2(n773), .Z(n775) );
  inv1 U695 ( .I(n956), .ZN(n687) );
  and2 U696 ( .A1(h2), .A2(f2), .Z(n617) );
  inv1 U697 ( .I(i3), .ZN(n431) );
  or2 U698 ( .A1(n616), .A2(n611), .Z(n695) );
  and2 U699 ( .A1(n970), .A2(n968), .Z(n726) );
  inv1 U700 ( .I(l2), .ZN(n924) );
  or2 U701 ( .A1(n852), .A2(n851), .Z(n863) );
  inv1 U702 ( .I(n850), .ZN(n852) );
  or2 U703 ( .A1(n846), .A2(n845), .Z(n847) );
  inv1 U704 ( .I(n651), .ZN(n865) );
  inv1 U705 ( .I(n903), .ZN(n922) );
  inv1 U706 ( .I(n363), .ZN(n928) );
  and2 U707 ( .A1(n890), .A2(n889), .Z(n891) );
  inv1 U708 ( .I(w2), .ZN(n729) );
  inv1 U709 ( .I(n790), .ZN(p4) );
  or2 U710 ( .A1(n815), .A2(n814), .Z(n816) );
  and2 U711 ( .A1(n825), .A2(n826), .Z(v4) );
  or2 U712 ( .A1(n1002), .A2(r2), .Z(n825) );
  inv1 U713 ( .I(n864), .ZN(n855) );
  inv1 U715 ( .I(n1002), .ZN(n1003) );
  inv1 U716 ( .I(r1), .ZN(n925) );
  and2 U717 ( .A1(n766), .A2(n947), .Z(n772) );
  and2 U718 ( .A1(n955), .A2(n767), .Z(n947) );
  and2f U719 ( .A1(n983), .A2(n763), .Z(n948) );
  inv1 U721 ( .I(d0), .ZN(n911) );
  and2f U722 ( .A1(n747), .A2(y3), .Z(n690) );
  or2 U723 ( .A1(n427), .A2(n952), .Z(n950) );
  and2 U724 ( .A1(n950), .A2(n951), .Z(n949) );
  inv1 U725 ( .I(n949), .ZN(n993) );
  or2 U726 ( .A1(n139), .A2(n304), .Z(n951) );
  or2 U727 ( .A1(n701), .A2(n139), .Z(n952) );
  inv1 U728 ( .I(n937), .ZN(n953) );
  buf0 U729 ( .I(n732), .Z(n954) );
  inv1 U730 ( .I(n932), .ZN(n955) );
  or2f U731 ( .A1(n997), .A2(z3), .Z(n956) );
  or2f U732 ( .A1(n958), .A2(n686), .Z(n957) );
  inv1f U733 ( .I(n979), .ZN(n937) );
  and2f U735 ( .A1(n768), .A2(n687), .Z(n958) );
  or2f U737 ( .A1(n651), .A2(n853), .Z(n854) );
  or2f U739 ( .A1(n509), .A2(n510), .Z(n184) );
  and2 U740 ( .A1(n400), .A2(n303), .Z(n409) );
  inv1 U742 ( .I(n303), .ZN(n410) );
  inv1 U743 ( .I(n467), .ZN(n774) );
  or2 U744 ( .A1(n938), .A2(n848), .Z(n960) );
  or2 U746 ( .A1(n845), .A2(n938), .Z(n961) );
  inv1f U747 ( .I(n997), .ZN(n998) );
  or2f U752 ( .A1(n700), .A2(n496), .Z(n903) );
  and2f U753 ( .A1(u2), .A2(n998), .Z(n870) );
  or2f U757 ( .A1(n781), .A2(n962), .Z(n790) );
  or2 U758 ( .A1(n780), .A2(n788), .Z(n962) );
  and2f U759 ( .A1(n964), .A2(n965), .Z(n963) );
  inv1f U760 ( .I(m), .ZN(n964) );
  inv1f U761 ( .I(d0), .ZN(n965) );
  or2f U762 ( .A1(n966), .A2(n981), .Z(n731) );
  or2f U763 ( .A1(n980), .A2(n729), .Z(n966) );
  and2 U764 ( .A1(n776), .A2(n775), .Z(n778) );
  and2 U765 ( .A1(n773), .A2(n776), .Z(n653) );
  inv1 U766 ( .I(n898), .ZN(n899) );
  and2f U767 ( .A1(n759), .A2(n690), .Z(n996) );
  and2f U768 ( .A1(n967), .A2(u2), .Z(n968) );
  inv1f U769 ( .I(n703), .ZN(n967) );
  and2 U770 ( .A1(n967), .A2(n970), .Z(n969) );
  or2f U771 ( .A1(s0), .A2(n971), .Z(n970) );
  and2f U772 ( .A1(n970), .A2(x2), .Z(n972) );
  and2f U773 ( .A1(n731), .A2(n760), .Z(n973) );
  inv1f U774 ( .I(n973), .ZN(n983) );
  or2f U775 ( .A1(h2), .A2(f2), .Z(n974) );
  inv1f U776 ( .I(n974), .ZN(n320) );
  inv1 U777 ( .I(h2), .ZN(n277) );
  inv1 U778 ( .I(f2), .ZN(n380) );
  or2f U779 ( .A1(n467), .A2(n925), .Z(n975) );
  inv1f U780 ( .I(n975), .ZN(n979) );
  and2 U781 ( .A1(y2), .A2(g3), .Z(n976) );
  or2 U782 ( .A1(n953), .A2(n978), .Z(n977) );
  or2 U784 ( .A1(p1), .A2(n320), .Z(n616) );
  and2f U785 ( .A1(n725), .A2(n982), .Z(n980) );
  and2f U786 ( .A1(n972), .A2(n968), .Z(n982) );
  or2f U787 ( .A1(n813), .A2(n948), .Z(n984) );
  inv1 U788 ( .I(s0), .ZN(n868) );
  and2f U791 ( .A1(n732), .A2(n987), .Z(n985) );
  or2f U792 ( .A1(n985), .A2(n986), .Z(n691) );
  and2 U793 ( .A1(n759), .A2(n729), .Z(n986) );
  and2 U794 ( .A1(x2), .A2(n759), .Z(n987) );
  inv1f U795 ( .I(n692), .ZN(n988) );
  or2f U797 ( .A1(n958), .A2(n686), .Z(n989) );
  or2 U798 ( .A1(n655), .A2(n916), .Z(n759) );
  inv1 U799 ( .I(n969), .ZN(n851) );
  or2f U800 ( .A1(n855), .A2(n990), .Z(n861) );
  or2 U802 ( .A1(n854), .A2(n858), .Z(n990) );
  and2f U803 ( .A1(n847), .A2(n993), .Z(n991) );
  or2f U809 ( .A1(n991), .A2(n992), .Z(n866) );
  and2 U810 ( .A1(n865), .A2(n938), .Z(n992) );
  and2f U811 ( .A1(n776), .A2(n775), .Z(n994) );
  or2f U812 ( .A1(n994), .A2(n995), .Z(n902) );
  or2 U813 ( .A1(n779), .A2(n777), .Z(n995) );
  and2f U814 ( .A1(n731), .A2(n996), .Z(n688) );
  inv1f U815 ( .I(n902), .ZN(n997) );
  and2f U816 ( .A1(n937), .A2(n976), .Z(n999) );
  or2f U817 ( .A1(n1001), .A2(n977), .Z(n1000) );
  inv1 U818 ( .I(n1000), .ZN(n684) );
  or2f U819 ( .A1(n772), .A2(n771), .Z(n1002) );
  or2 U820 ( .A1(n998), .A2(n901), .Z(n906) );
  and2 U822 ( .A1(a), .A2(f0), .Z(n777) );
  or2 U823 ( .A1(z2), .A2(a3), .Z(n701) );
  inv1 U824 ( .I(r2), .ZN(n779) );
  or2 U825 ( .A1(n886), .A2(n699), .Z(n938) );
  inv1 U826 ( .I(a2), .ZN(n699) );
  and2 U827 ( .A1(s0), .A2(n751), .Z(n752) );
  inv1 U828 ( .I(n459), .ZN(n751) );
  and2 U829 ( .A1(b2), .A2(n288), .Z(n459) );
  inv1 U830 ( .I(n458), .ZN(n753) );
  or2 U831 ( .A1(t1), .A2(n706), .Z(n322) );
  inv1 U832 ( .I(t2), .ZN(n706) );
  or2 U833 ( .A1(n266), .A2(o0), .Z(n261) );
  and2 U834 ( .A1(h2), .A2(n267), .Z(n266) );
  or2 U835 ( .A1(e3), .A2(n762), .Z(n763) );
  or2 U843 ( .A1(f3), .A2(n757), .Z(n761) );
  and2 U844 ( .A1(n929), .A2(m3), .Z(n757) );
  or2 U845 ( .A1(n927), .A2(n222), .Z(n828) );
  and2 U846 ( .A1(n224), .A2(n), .Z(n222) );
  and2 U847 ( .A1(n656), .A2(n226), .Z(n224) );
  inv1 U848 ( .I(n828), .ZN(n829) );
  or2 U849 ( .A1(n738), .A2(l3), .Z(n845) );
  inv1 U850 ( .I(y), .ZN(n579) );
  inv1 U853 ( .I(n498), .ZN(n856) );
  and2 U854 ( .A1(l0), .A2(m0), .Z(n498) );
  or2 U855 ( .A1(n130), .A2(n499), .Z(n496) );
  inv1 U857 ( .I(k0), .ZN(n499) );
  or2 U860 ( .A1(h3), .A2(n431), .Z(n170) );
  or2 U861 ( .A1(n400), .A2(n929), .Z(n304) );
  inv1 U862 ( .I(o), .ZN(n171) );
  or2 U863 ( .A1(n930), .A2(n500), .Z(n244) );
  or2 U865 ( .A1(n501), .A2(n502), .Z(n500) );
  inv1 U866 ( .I(n184), .ZN(n930) );
  and2 U867 ( .A1(z0), .A2(w0), .Z(n502) );
  inv1 U868 ( .I(q), .ZN(n169) );
  inv1 U872 ( .I(n560), .ZN(n555) );
  and2 U873 ( .A1(w2), .A2(n770), .Z(n771) );
  or2 U874 ( .A1(n916), .A2(n769), .Z(n770) );
  and2 U875 ( .A1(n655), .A2(n915), .Z(n769) );
  inv1 U876 ( .I(n1), .ZN(n748) );
  inv1 U879 ( .I(v2), .ZN(n893) );
  inv1 U881 ( .I(n578), .ZN(n577) );
  and2 U882 ( .A1(n579), .A2(x), .Z(n578) );
  inv1 U883 ( .I(n745), .ZN(n746) );
  or2 U884 ( .A1(n744), .A2(n743), .Z(n745) );
  and2 U885 ( .A1(n526), .A2(n742), .Z(n744) );
  and2 U886 ( .A1(n564), .A2(n565), .Z(n415) );
  and2 U888 ( .A1(x1), .A2(r0), .Z(n565) );
  and2 U889 ( .A1(m2), .A2(n566), .Z(n564) );
  and2 U890 ( .A1(n176), .A2(n555), .Z(n566) );
  and2 U891 ( .A1(n417), .A2(n418), .Z(n416) );
  or2 U892 ( .A1(n419), .A2(n420), .Z(n418) );
  inv1 U893 ( .I(w1), .ZN(n175) );
  inv1 U895 ( .I(n322), .ZN(n780) );
  and2 U896 ( .A1(n786), .A2(n785), .Z(n787) );
  and2 U897 ( .A1(n974), .A2(n783), .Z(n785) );
  inv1 U899 ( .I(n375), .ZN(n786) );
  or2 U900 ( .A1(n782), .A2(n366), .Z(n783) );
  inv1 U904 ( .I(n321), .ZN(n319) );
  or2 U905 ( .A1(n322), .A2(a), .Z(n321) );
  and2 U906 ( .A1(n262), .A2(n263), .Z(n259) );
  or2 U907 ( .A1(g2), .A2(n264), .Z(n263) );
  and2 U908 ( .A1(n265), .A2(n261), .Z(n262) );
  or2 U909 ( .A1(n268), .A2(n269), .Z(n265) );
  and2 U910 ( .A1(n261), .A2(n924), .Z(n260) );
  or2 U912 ( .A1(n274), .A2(n275), .Z(n273) );
  and2 U913 ( .A1(n283), .A2(n284), .Z(n274) );
  and2 U915 ( .A1(n268), .A2(n276), .Z(n275) );
  and2 U916 ( .A1(n285), .A2(n286), .Z(n284) );
  inv1 U917 ( .I(a), .ZN(n927) );
  inv1 U918 ( .I(n653), .ZN(n931) );
  or2 U919 ( .A1(n828), .A2(n2), .Z(n821) );
  inv1 U924 ( .I(n820), .ZN(n823) );
  or2 U926 ( .A1(n828), .A2(n827), .Z(n836) );
  inv1 U927 ( .I(b), .ZN(n827) );
  or2 U928 ( .A1(n829), .A2(b), .Z(n830) );
  or2 U932 ( .A1(n834), .A2(c), .Z(n838) );
  inv1 U933 ( .I(n836), .ZN(n834) );
  or2 U934 ( .A1(n836), .A2(n835), .Z(n837) );
  inv1 U935 ( .I(c), .ZN(n835) );
  inv1 U936 ( .I(n481), .ZN(n622) );
  and2 U937 ( .A1(c1), .A2(d1), .Z(n481) );
  inv1 U938 ( .I(e1), .ZN(n603) );
  and2 U939 ( .A1(n603), .A2(l2), .Z(n568) );
  and2 U940 ( .A1(n491), .A2(n522), .Z(n550) );
  inv1 U941 ( .I(d1), .ZN(n522) );
  inv1 U942 ( .I(c1), .ZN(n491) );
  and2 U943 ( .A1(n601), .A2(l2), .Z(n490) );
  or2 U944 ( .A1(n602), .A2(n169), .Z(n601) );
  or2 U945 ( .A1(n420), .A2(p), .Z(n602) );
  inv1 U946 ( .I(n441), .ZN(n226) );
  and2 U947 ( .A1(n442), .A2(f), .Z(n441) );
  and2 U948 ( .A1(e), .A2(d), .Z(n442) );
  and2 U949 ( .A1(n380), .A2(g2), .Z(n404) );
  and2 U950 ( .A1(l2), .A2(g2), .Z(n366) );
  and2 U951 ( .A1(f2), .A2(l2), .Z(n367) );
  or2 U952 ( .A1(n856), .A2(n496), .Z(n857) );
  inv1 U953 ( .I(o3), .ZN(n945) );
  inv1 U954 ( .I(n938), .ZN(n923) );
  or2 U955 ( .A1(n701), .A2(h0), .Z(n843) );
  or2 U956 ( .A1(n938), .A2(n868), .Z(n869) );
  and2 U957 ( .A1(n173), .A2(n174), .Z(n172) );
  and2 U958 ( .A1(n175), .A2(n176), .Z(n174) );
  or2 U959 ( .A1(n164), .A2(n165), .Z(n163) );
  and2 U960 ( .A1(n167), .A2(n166), .Z(n164) );
  and2 U961 ( .A1(n166), .A2(p2), .Z(n165) );
  and2 U962 ( .A1(n170), .A2(n171), .Z(n167) );
  or2 U963 ( .A1(n845), .A2(n486), .Z(n936) );
  or2 U964 ( .A1(g0), .A2(n971), .Z(n486) );
  or2 U965 ( .A1(n740), .A2(n739), .Z(n848) );
  or2 U966 ( .A1(n738), .A2(n737), .Z(n739) );
  or2 U967 ( .A1(l2), .A2(n184), .Z(n740) );
  inv1 U968 ( .I(g0), .ZN(n737) );
  and2 U969 ( .A1(n244), .A2(j2), .Z(n130) );
  inv1 U970 ( .I(n697), .ZN(n128) );
  or2 U971 ( .A1(n696), .A2(n738), .Z(n697) );
  inv1 U972 ( .I(n520), .ZN(n696) );
  and2 U973 ( .A1(n971), .A2(n3), .Z(n520) );
  inv1 U974 ( .I(n649), .ZN(n650) );
  or2 U975 ( .A1(x), .A2(n579), .Z(n649) );
  inv1 U976 ( .I(y1), .ZN(n176) );
  or2 U977 ( .A1(n944), .A2(q2), .Z(n584) );
  inv1 U978 ( .I(p2), .ZN(n944) );
  inv1 U979 ( .I(p0), .ZN(n548) );
  inv1 U980 ( .I(n544), .ZN(n542) );
  or2 U981 ( .A1(n563), .A2(n415), .Z(n544) );
  and2 U982 ( .A1(n567), .A2(n560), .Z(n563) );
  and2 U983 ( .A1(p), .A2(n558), .Z(n567) );
  or2 U984 ( .A1(n545), .A2(n546), .Z(n543) );
  and2 U985 ( .A1(q0), .A2(n548), .Z(n545) );
  inv1 U986 ( .I(n547), .ZN(n546) );
  or2 U987 ( .A1(n548), .A2(q0), .Z(n547) );
  or2 U988 ( .A1(n495), .A2(n856), .Z(n700) );
  and2 U989 ( .A1(n517), .A2(n518), .Z(n495) );
  or2 U990 ( .A1(n924), .A2(n555), .Z(n488) );
  and2 U991 ( .A1(m2), .A2(n170), .Z(n480) );
  inv1 U992 ( .I(k2), .ZN(n479) );
  and2 U993 ( .A1(n482), .A2(n479), .Z(n943) );
  inv1 U994 ( .I(m0), .ZN(n482) );
  inv1 U995 ( .I(n936), .ZN(n920) );
  and2 U996 ( .A1(n918), .A2(n424), .Z(n408) );
  inv1 U997 ( .I(n843), .ZN(n918) );
  and2 U998 ( .A1(n399), .A2(t0), .Z(n424) );
  and2 U999 ( .A1(n431), .A2(h3), .Z(n400) );
  inv1 U1000 ( .I(n304), .ZN(n390) );
  and2 U1001 ( .A1(n919), .A2(n399), .Z(n391) );
  inv1 U1002 ( .I(n701), .ZN(n919) );
  inv1 U1003 ( .I(o0), .ZN(n241) );
  or2 U1004 ( .A1(n171), .A2(n208), .Z(n140) );
  or2 U1005 ( .A1(n209), .A2(n924), .Z(n208) );
  and2 U1006 ( .A1(j2), .A2(n243), .Z(n206) );
  inv1 U1007 ( .I(n244), .ZN(n243) );
  or2 U1008 ( .A1(n515), .A2(n516), .Z(n509) );
  or2 U1009 ( .A1(n511), .A2(n512), .Z(n510) );
  and2 U1010 ( .A1(y0), .A2(n508), .Z(n515) );
  or2 U1011 ( .A1(n288), .A2(n467), .Z(n596) );
  and2 U1012 ( .A1(o1), .A2(n608), .Z(n599) );
  inv1 U1013 ( .I(y3), .ZN(n608) );
  or2 U1014 ( .A1(n595), .A2(n924), .Z(n593) );
  and2 U1015 ( .A1(m1), .A2(n596), .Z(n595) );
  or2 U1016 ( .A1(n169), .A2(n572), .Z(n594) );
  or2 U1017 ( .A1(n169), .A2(n488), .Z(n598) );
  or2 U1018 ( .A1(n599), .A2(i1), .Z(n597) );
  or2 U1019 ( .A1(l3), .A2(s), .Z(n458) );
  or2 U1020 ( .A1(p2), .A2(q2), .Z(n572) );
  inv1 U1021 ( .I(k1), .ZN(n539) );
  inv1 U1022 ( .I(n535), .ZN(n533) );
  or2 U1023 ( .A1(n553), .A2(n554), .Z(n535) );
  and2 U1024 ( .A1(n559), .A2(q), .Z(n553) );
  and2 U1025 ( .A1(n417), .A2(n555), .Z(n554) );
  and2 U1026 ( .A1(n560), .A2(n558), .Z(n559) );
  or2 U1027 ( .A1(n536), .A2(n537), .Z(n534) );
  and2 U1028 ( .A1(l1), .A2(n539), .Z(n536) );
  inv1 U1029 ( .I(n538), .ZN(n537) );
  or2 U1030 ( .A1(n539), .A2(l1), .Z(n538) );
  and2 U1031 ( .A1(i1), .A2(n581), .Z(n940) );
  and2 U1032 ( .A1(y3), .A2(e4), .Z(n581) );
  and2 U1033 ( .A1(y1), .A2(n556), .Z(n417) );
  inv1 U1034 ( .I(n557), .ZN(n556) );
  or2 U1035 ( .A1(x1), .A2(n558), .Z(n557) );
  inv1 U1036 ( .I(l3), .ZN(n880) );
  or2 U1037 ( .A1(n698), .A2(n3), .Z(n885) );
  or2 U1038 ( .A1(t3), .A2(o3), .Z(n698) );
  or2 U1039 ( .A1(n749), .A2(n748), .Z(n887) );
  and2 U1040 ( .A1(n691), .A2(n747), .Z(n749) );
  inv1 U1041 ( .I(n885), .ZN(n886) );
  inv1 U1042 ( .I(s1), .ZN(n288) );
  and2 U1043 ( .A1(n925), .A2(s1), .Z(n656) );
  or2 U1044 ( .A1(k3), .A2(n137), .Z(n136) );
  inv1 U1045 ( .I(p3), .ZN(n137) );
  inv1 U1046 ( .I(n954), .ZN(n915) );
  inv1 U1047 ( .I(n655), .ZN(n939) );
  and2 U1048 ( .A1(x0), .A2(n159), .Z(n506) );
  and2 U1049 ( .A1(n171), .A2(n279), .Z(n267) );
  inv1 U1050 ( .I(n209), .ZN(n279) );
  inv1 U1051 ( .I(f1), .ZN(n272) );
  and2 U1052 ( .A1(n291), .A2(n292), .Z(n271) );
  inv1 U1053 ( .I(g1), .ZN(n291) );
  inv1 U1054 ( .I(h1), .ZN(n292) );
  and2 U1055 ( .A1(v1), .A2(b2), .Z(n758) );
  or2 U1056 ( .A1(n436), .A2(n437), .Z(n435) );
  and2 U1057 ( .A1(o0), .A2(l2), .Z(n436) );
  inv1 U1058 ( .I(n438), .ZN(n437) );
  or2 U1059 ( .A1(d3), .A2(b3), .Z(n438) );
  inv1 U1060 ( .I(c3), .ZN(n434) );
  inv1 U1061 ( .I(n170), .ZN(n929) );
  and2 U1062 ( .A1(n503), .A2(n504), .Z(n501) );
  and2 U1063 ( .A1(n508), .A2(n158), .Z(n503) );
  or2 U1064 ( .A1(n505), .A2(n506), .Z(n504) );
  and2 U1065 ( .A1(y0), .A2(n507), .Z(n505) );
  or2 U1066 ( .A1(s1), .A2(n925), .Z(n613) );
  and2 U1067 ( .A1(u2), .A2(n754), .Z(n755) );
  or2 U1068 ( .A1(n753), .A2(n752), .Z(n754) );
  or2 U1069 ( .A1(n741), .A2(t), .Z(n742) );
  or2 U1070 ( .A1(n971), .A2(n527), .Z(n526) );
  or2 U1071 ( .A1(s0), .A2(g0), .Z(n527) );
  inv1 U1072 ( .I(u2), .ZN(n743) );
  inv1 U1073 ( .I(z1), .ZN(n782) );
  and2 U1074 ( .A1(n376), .A2(n377), .Z(n375) );
  or2 U1075 ( .A1(n380), .A2(n277), .Z(n376) );
  or2 U1076 ( .A1(n378), .A2(z1), .Z(n377) );
  inv1 U1077 ( .I(n379), .ZN(n378) );
  and2 U1078 ( .A1(n270), .A2(n271), .Z(n269) );
  and2 U1079 ( .A1(g2), .A2(n272), .Z(n270) );
  and2 U1080 ( .A1(n925), .A2(n288), .Z(n285) );
  inv1 U1081 ( .I(q1), .ZN(n286) );
  or2 U1082 ( .A1(n277), .A2(n278), .Z(n276) );
  or2 U1083 ( .A1(o0), .A2(n267), .Z(n278) );
  inv1 U1084 ( .I(n280), .ZN(n268) );
  or2 U1085 ( .A1(n281), .A2(n282), .Z(n280) );
  or2 U1086 ( .A1(s1), .A2(r1), .Z(n281) );
  or2 U1087 ( .A1(q1), .A2(g2), .Z(n282) );
  and2 U1088 ( .A1(n289), .A2(n277), .Z(n283) );
  or2 U1089 ( .A1(n290), .A2(n924), .Z(n289) );
  and2 U1090 ( .A1(n271), .A2(n272), .Z(n290) );
  or2 U1091 ( .A1(n969), .A2(n743), .Z(n773) );
  inv1 U1092 ( .I(c2), .ZN(n735) );
  inv1 U1093 ( .I(o2), .ZN(n803) );
  inv1 U1094 ( .I(n2), .ZN(n804) );
  inv1 U1095 ( .I(n), .ZN(n420) );
  and2 U1096 ( .A1(u2), .A2(n843), .Z(n844) );
  and2 U1097 ( .A1(p), .A2(n168), .Z(n166) );
  and2 U1098 ( .A1(n169), .A2(l2), .Z(n168) );
  inv1 U1099 ( .I(t0), .ZN(n738) );
  or2 U1100 ( .A1(n128), .A2(n938), .Z(n518) );
  inv1 U1101 ( .I(j0), .ZN(n517) );
  inv1 U1102 ( .I(m3), .ZN(n395) );
  or2 U1103 ( .A1(n432), .A2(n433), .Z(n425) );
  and2 U1104 ( .A1(n439), .A2(o0), .Z(n432) );
  and2 U1105 ( .A1(n434), .A2(n435), .Z(n433) );
  and2 U1106 ( .A1(d3), .A2(l2), .Z(n439) );
  or2 U1107 ( .A1(n395), .A2(n396), .Z(n394) );
  or2 U1108 ( .A1(n979), .A2(n390), .Z(n396) );
  or2 U1109 ( .A1(n430), .A2(n431), .Z(n393) );
  inv1 U1110 ( .I(h3), .ZN(n430) );
  inv1 U1111 ( .I(n425), .ZN(n399) );
  and2 U1112 ( .A1(a3), .A2(n851), .Z(n704) );
  inv1 U1113 ( .I(u), .ZN(n354) );
  or2 U1114 ( .A1(n937), .A2(z2), .Z(n360) );
  or2 U1115 ( .A1(p), .A2(q), .Z(n209) );
  or2 U1116 ( .A1(n513), .A2(n514), .Z(n512) );
  and2 U1117 ( .A1(z0), .A2(n507), .Z(n513) );
  and2 U1118 ( .A1(x0), .A2(n158), .Z(n514) );
  inv1 U1119 ( .I(u1), .ZN(n511) );
  and2 U1120 ( .A1(w0), .A2(n159), .Z(n516) );
  inv1 U1121 ( .I(y0), .ZN(n159) );
  inv1 U1122 ( .I(z0), .ZN(n158) );
  and2 U1123 ( .A1(p2), .A2(q2), .Z(n560) );
  inv1 U1124 ( .I(m2), .ZN(n558) );
  inv1 U1125 ( .I(z3), .ZN(n767) );
  and2 U1126 ( .A1(b2), .A2(n656), .Z(n747) );
  inv1 U1127 ( .I(x0), .ZN(n507) );
  inv1 U1128 ( .I(w0), .ZN(n508) );
  and2 U1129 ( .A1(y2), .A2(n984), .Z(n799) );
  and2 U1130 ( .A1(n796), .A2(n793), .Z(n801) );
  or2 U1131 ( .A1(n792), .A2(n235), .Z(n793) );
  and2 U1132 ( .A1(v), .A2(s0), .Z(n235) );
  inv1 U1133 ( .I(n807), .ZN(n808) );
  and2 U1134 ( .A1(n806), .A2(n805), .Z(n807) );
  or2 U1135 ( .A1(n829), .A2(n804), .Z(n805) );
  or2 U1136 ( .A1(n821), .A2(n803), .Z(n806) );
  and2 U1137 ( .A1(n813), .A2(n812), .Z(n815) );
  and2 U1138 ( .A1(y2), .A2(n811), .Z(n812) );
  and2 U1139 ( .A1(o2), .A2(n821), .Z(n817) );
  and2 U1140 ( .A1(e1), .A2(n481), .Z(n419) );
  or2 U1141 ( .A1(n355), .A2(n356), .Z(n350) );
  and2 U1142 ( .A1(n868), .A2(n705), .Z(n356) );
  and2 U1143 ( .A1(n360), .A2(n704), .Z(n355) );
  and2 U1144 ( .A1(i0), .A2(n971), .Z(n705) );
  or2 U1145 ( .A1(n352), .A2(n304), .Z(n351) );
  and2 U1146 ( .A1(n353), .A2(v), .Z(n352) );
  and2 U1147 ( .A1(s0), .A2(n354), .Z(n353) );
  and2 U1148 ( .A1(n363), .A2(n360), .Z(n362) );
  and2 U1149 ( .A1(n158), .A2(n159), .Z(n941) );
  inv1 U1150 ( .I(y2), .ZN(n889) );
  or2 U1151 ( .A1(n904), .A2(n922), .Z(n905) );
  and2 U1152 ( .A1(i1), .A2(e4), .Z(n904) );
  or2 U1153 ( .A1(n734), .A2(d4), .Z(n249) );
  or2 U1154 ( .A1(n913), .A2(n932), .Z(n734) );
  inv1 U1155 ( .I(n733), .ZN(n913) );
  or2 U1156 ( .A1(n915), .A2(n939), .Z(n733) );
  and2 U1157 ( .A1(n507), .A2(n508), .Z(n942) );
  inv1 U1158 ( .I(x2), .ZN(n916) );
  and2 U1159 ( .A1(j1), .A2(n578), .Z(n575) );
  and2 U1160 ( .A1(e0), .A2(n577), .Z(n576) );
  and2 U1161 ( .A1(k1), .A2(y1), .Z(n569) );
  and2 U1162 ( .A1(p0), .A2(n176), .Z(n570) );
  and2 U1163 ( .A1(n655), .A2(n175), .Z(n413) );
  or2 U1164 ( .A1(n415), .A2(n416), .Z(n414) );
  or2 U1165 ( .A1(n787), .A2(a), .Z(n788) );
  and2 U1166 ( .A1(a1), .A2(t2), .Z(n318) );
  and2 U1167 ( .A1(n319), .A2(n320), .Z(n317) );
  and2 U1168 ( .A1(a), .A2(n273), .Z(n257) );
  or2 U1169 ( .A1(n259), .A2(n260), .Z(n258) );
  or2 U1170 ( .A1(n736), .A2(f0), .Z(n246) );
  and2 U1171 ( .A1(n931), .A2(n774), .Z(n736) );
  and2 U1172 ( .A1(n823), .A2(n822), .Z(n826) );
  or2 U1173 ( .A1(n821), .A2(o2), .Z(n822) );
  and2 U1174 ( .A1(n836), .A2(n830), .Z(n831) );
  and2 U1175 ( .A1(n838), .A2(n837), .Z(n839) );
  and2 U1176 ( .A1(v0), .A2(n133), .Z(n132) );
  inv1 U1177 ( .I(x3), .ZN(n133) );
  and2 U1178 ( .A1(d1), .A2(n491), .Z(n626) );
  and2 U1179 ( .A1(c1), .A2(n522), .Z(n627) );
  and2 U1180 ( .A1(n481), .A2(n603), .Z(n621) );
  and2 U1181 ( .A1(e1), .A2(n622), .Z(n620) );
  and2 U1182 ( .A1(n550), .A2(n568), .Z(n600) );
  and2 U1183 ( .A1(n568), .A2(n522), .Z(n585) );
  and2 U1184 ( .A1(n568), .A2(n491), .Z(n574) );
  and2 U1185 ( .A1(n550), .A2(l2), .Z(n549) );
  and2 U1186 ( .A1(l2), .A2(n522), .Z(n521) );
  and2 U1187 ( .A1(l2), .A2(n491), .Z(n489) );
  or2 U1188 ( .A1(n656), .A2(b1), .Z(n440) );
  and2 U1189 ( .A1(n412), .A2(n404), .Z(n411) );
  and2 U1190 ( .A1(h2), .A2(n924), .Z(n412) );
  or2 U1191 ( .A1(n403), .A2(n277), .Z(n402) );
  or2 U1192 ( .A1(n404), .A2(l2), .Z(n403) );
  and2 U1193 ( .A1(n277), .A2(n924), .Z(n364) );
  or2 U1194 ( .A1(n366), .A2(n367), .Z(n365) );
  or2 U1195 ( .A1(n923), .A2(j0), .Z(n860) );
  or2 U1196 ( .A1(n857), .A2(n128), .Z(n858) );
  and2 U1197 ( .A1(n863), .A2(n862), .Z(n867) );
  and2 U1198 ( .A1(n936), .A2(n922), .Z(n862) );
  and2 U1199 ( .A1(n923), .A2(n945), .Z(n242) );
  and2 U1200 ( .A1(k0), .A2(n212), .Z(n211) );
  or2 U1201 ( .A1(n938), .A2(n843), .Z(n212) );
  inv1 U1202 ( .I(n873), .ZN(n874) );
  or2 U1203 ( .A1(n162), .A2(n163), .Z(n160) );
  or2 U1204 ( .A1(m0), .A2(n172), .Z(n162) );
  and2 U1205 ( .A1(k2), .A2(n140), .Z(n138) );
  inv1 U1206 ( .I(n848), .ZN(n139) );
  and2 U1207 ( .A1(n131), .A2(l3), .Z(n129) );
  and2 U1208 ( .A1(g0), .A2(t0), .Z(n131) );
  or2 U1209 ( .A1(k2), .A2(i2), .Z(n126) );
  or2 U1210 ( .A1(n128), .A2(n932), .Z(n876) );
  and2 U1211 ( .A1(n0), .A2(n649), .Z(n648) );
  and2 U1212 ( .A1(n650), .A2(e0), .Z(n647) );
  or2 U1213 ( .A1(m1), .A2(n625), .Z(n624) );
  or2 U1214 ( .A1(r0), .A2(q2), .Z(n625) );
  and2 U1215 ( .A1(w1), .A2(x1), .Z(n618) );
  and2 U1216 ( .A1(m2), .A2(n176), .Z(n619) );
  and2 U1217 ( .A1(q2), .A2(n944), .Z(n582) );
  inv1 U1218 ( .I(n584), .ZN(n583) );
  or2 U1219 ( .A1(r0), .A2(n572), .Z(n573) );
  and2 U1220 ( .A1(n544), .A2(n548), .Z(n562) );
  and2 U1221 ( .A1(v3), .A2(n542), .Z(n561) );
  and2 U1222 ( .A1(n543), .A2(n544), .Z(n540) );
  and2 U1223 ( .A1(w3), .A2(n542), .Z(n541) );
  and2 U1224 ( .A1(n487), .A2(r0), .Z(n484) );
  and2 U1225 ( .A1(n488), .A2(n937), .Z(n487) );
  and2 U1226 ( .A1(n478), .A2(n479), .Z(n477) );
  or2 U1227 ( .A1(n480), .A2(p2), .Z(n478) );
  or2 U1228 ( .A1(n408), .A2(n920), .Z(n423) );
  and2 U1229 ( .A1(n410), .A2(h3), .Z(n422) );
  or2 U1230 ( .A1(n406), .A2(n407), .Z(n6) );
  and2 U1231 ( .A1(n410), .A2(i3), .Z(n406) );
  or2 U1232 ( .A1(n408), .A2(n409), .Z(n407) );
  or2 U1233 ( .A1(n878), .A2(n387), .Z(o6) );
  and2 U1234 ( .A1(n928), .A2(n969), .Z(n878) );
  and2 U1235 ( .A1(z2), .A2(n389), .Z(n387) );
  or2 U1236 ( .A1(n346), .A2(n347), .Z(p6) );
  and2 U1237 ( .A1(n928), .A2(n349), .Z(n347) );
  and2 U1238 ( .A1(n362), .A2(a3), .Z(n346) );
  or2 U1239 ( .A1(n350), .A2(n351), .Z(n349) );
  and2 U1240 ( .A1(n251), .A2(n241), .Z(n250) );
  or2 U1241 ( .A1(b3), .A2(n937), .Z(n251) );
  and2 U1242 ( .A1(c3), .A2(o0), .Z(n240) );
  and2 U1243 ( .A1(d3), .A2(n241), .Z(n239) );
  inv1 U1244 ( .I(n207), .ZN(n205) );
  or2 U1245 ( .A1(n140), .A2(k2), .Z(n207) );
  and2 U1246 ( .A1(t0), .A2(n184), .Z(n183) );
  or2 U1247 ( .A1(n599), .A2(m1), .Z(n607) );
  and2 U1248 ( .A1(n596), .A2(n598), .Z(n606) );
  and2 U1249 ( .A1(n597), .A2(n598), .Z(n591) );
  or2 U1250 ( .A1(n593), .A2(n594), .Z(n592) );
  and2 U1251 ( .A1(n940), .A2(n458), .Z(n580) );
  or2 U1252 ( .A1(m1), .A2(n572), .Z(n571) );
  and2 U1253 ( .A1(n535), .A2(n539), .Z(n552) );
  and2 U1254 ( .A1(q3), .A2(n533), .Z(n551) );
  and2 U1255 ( .A1(n534), .A2(n535), .Z(n531) );
  and2 U1256 ( .A1(r3), .A2(n533), .Z(n532) );
  and2 U1257 ( .A1(s), .A2(n880), .Z(n881) );
  and2 U1258 ( .A1(n885), .A2(n884), .Z(m7) );
  or2 U1259 ( .A1(n888), .A2(n895), .Z(o7) );
  and2 U1260 ( .A1(u0), .A2(s2), .Z(n135) );
  and2 U1261 ( .A1(r), .A2(n136), .Z(n134) );
  and2 U1262 ( .A1(m), .A2(d0), .Z(n124) );
  and2 U1263 ( .A1(k), .A2(n911), .Z(n912) );
  and2 U1264 ( .A1(n623), .A2(n655), .Z(n914) );
  and2 U1265 ( .A1(x2), .A2(n729), .Z(n623) );
  inv1 U1266 ( .I(a4), .ZN(n605) );
  and2 U1267 ( .A1(w2), .A2(n939), .Z(n604) );
  or2 U1268 ( .A1(n575), .A2(n576), .Z(f4) );
  or2 U1269 ( .A1(n569), .A2(n570), .Z(g4) );
  or2 U1270 ( .A1(n413), .A2(n414), .Z(n4) );
  and2 U1271 ( .A1(w1), .A2(n655), .Z(o4) );
  or2 U1272 ( .A1(n317), .A2(n318), .Z(q4) );
  or2 U1273 ( .A1(n257), .A2(n258), .Z(r4) );
  and2 U1274 ( .A1(n246), .A2(n927), .Z(s4) );
  or2 U1275 ( .A1(n132), .A2(a), .Z(y4) );
  and2 U1276 ( .A1(v0), .A2(b4), .Z(z4) );
  or2 U1277 ( .A1(n626), .A2(n627), .Z(b5) );
  or2 U1278 ( .A1(n620), .A2(n621), .Z(c5) );
  or2 U1279 ( .A1(n600), .A2(n490), .Z(d5) );
  or2 U1280 ( .A1(n585), .A2(n490), .Z(e5) );
  or2 U1281 ( .A1(n574), .A2(n490), .Z(f5) );
  or2 U1282 ( .A1(n568), .A2(n490), .Z(g5) );
  or2 U1283 ( .A1(n549), .A2(n490), .Z(h5) );
  or2 U1284 ( .A1(n521), .A2(n490), .Z(i5) );
  or2 U1285 ( .A1(n489), .A2(n490), .Z(j5) );
  and2 U1286 ( .A1(n419), .A2(n), .Z(l5) );
  and2 U1287 ( .A1(n440), .A2(n226), .Z(m5) );
  or2 U1288 ( .A1(n411), .A2(a), .Z(n5) );
  inv1 U1289 ( .I(n402), .ZN(o5) );
  or2 U1290 ( .A1(n364), .A2(n365), .Z(p5) );
  or2 U1291 ( .A1(n242), .A2(n206), .Z(s5) );
  or2 U1292 ( .A1(n211), .A2(l2), .Z(t5) );
  and2 U1293 ( .A1(n160), .A2(n936), .Z(v5) );
  and2 U1294 ( .A1(n922), .A2(n3), .Z(w5) );
  or2 U1295 ( .A1(n138), .A2(n139), .Z(x5) );
  or2 U1296 ( .A1(n129), .A2(n130), .Z(y5) );
  or2 U1297 ( .A1(n876), .A2(n126), .Z(z5) );
  or2 U1298 ( .A1(n647), .A2(n648), .Z(a6) );
  and2 U1299 ( .A1(m2), .A2(n624), .Z(b6) );
  and2 U1300 ( .A1(n618), .A2(n619), .Z(c6) );
  or2 U1301 ( .A1(n582), .A2(n583), .Z(e6) );
  and2 U1302 ( .A1(m2), .A2(n573), .Z(f6) );
  or2 U1303 ( .A1(n561), .A2(n562), .Z(g6) );
  or2 U1304 ( .A1(n540), .A2(n541), .Z(h6) );
  and2 U1305 ( .A1(n922), .A2(l3), .Z(i6) );
  or2 U1306 ( .A1(n484), .A2(n920), .Z(j6) );
  or2 U1307 ( .A1(n477), .A2(n943), .Z(l6) );
  or2 U1308 ( .A1(n422), .A2(n423), .Z(m6) );
  and2 U1309 ( .A1(b3), .A2(n241), .Z(q6) );
  and2 U1310 ( .A1(n250), .A2(c3), .Z(r6) );
  or2 U1311 ( .A1(n239), .A2(n240), .Z(s6) );
  or2 U1312 ( .A1(n205), .A2(n206), .Z(t6) );
  and2 U1313 ( .A1(n183), .A2(g0), .Z(u6) );
  and2 U1314 ( .A1(n606), .A2(n607), .Z(c7) );
  and2 U1315 ( .A1(n591), .A2(n592), .Z(d7) );
  and2 U1316 ( .A1(n580), .A2(z3), .Z(e7) );
  and2 U1317 ( .A1(m2), .A2(n571), .Z(f7) );
  or2 U1318 ( .A1(n551), .A2(n552), .Z(g7) );
  or2 U1319 ( .A1(n531), .A2(n532), .Z(h7) );
  inv1 U1320 ( .I(n879), .ZN(j7) );
  or2 U1321 ( .A1(n417), .A2(i1), .Z(k7) );
  and2 U1322 ( .A1(n249), .A2(n288), .Z(q7) );
  and2 U1323 ( .A1(n656), .A2(n249), .Z(r7) );
  or2 U1324 ( .A1(n134), .A2(n135), .Z(x7) );
  and2 U1325 ( .A1(p3), .A2(j3), .Z(y7) );
  or2 U1326 ( .A1(n912), .A2(n124), .Z(z7) );
  or2 U1327 ( .A1(n913), .A2(c4), .Z(a8) );
  and2 U1328 ( .A1(n915), .A2(n914), .Z(b8) );
  or2 U1329 ( .A1(n604), .A2(n605), .Z(c8) );
  and2 U1330 ( .A1(n729), .A2(n917), .Z(h8) );
endmodule

