
module term1 ( i0, h0, g0, f0, e0, d0, c0, a0, z, y, x, w, v, u, t, s, r, q, p, 
        o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, s0, r0, q0, p0, o0, n0, 
        m0, l0, k0, j0 );
  input i0, h0, g0, f0, e0, d0, c0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n,
         m, l, k, j, i, h, g, f, e, d, c, b, a;
  output s0, r0, q0, p0, o0, n0, m0, l0, k0, j0;
  wire   n304, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n305, n306, n307, n308, n309, n310, n311;

  or2f U4 ( .A1(n53), .A2(n52), .Z(n51) );
  and2f U5 ( .A1(n54), .A2(p), .Z(n53) );
  and2f U6 ( .A1(n55), .A2(n56), .Z(n54) );
  or2f U7 ( .A1(n57), .A2(n58), .Z(n55) );
  or2f U8 ( .A1(n59), .A2(n60), .Z(n58) );
  and2f U18 ( .A1(n74), .A2(n73), .Z(n59) );
  and2f U19 ( .A1(n75), .A2(n76), .Z(n74) );
  and2f U21 ( .A1(n77), .A2(n65), .Z(n75) );
  or2f U22 ( .A1(n78), .A2(n79), .Z(n77) );
  or2f U23 ( .A1(n311), .A2(n81), .Z(n79) );
  and2f U24 ( .A1(n82), .A2(n83), .Z(n73) );
  or2f U36 ( .A1(n98), .A2(n99), .Z(n97) );
  or2f U37 ( .A1(n100), .A2(n101), .Z(n99) );
  or2f U56 ( .A1(n118), .A2(n121), .Z(n84) );
  and2f U58 ( .A1(n66), .A2(n78), .Z(n118) );
  and2f U66 ( .A1(n138), .A2(n139), .Z(n80) );
  or2f U68 ( .A1(n141), .A2(n131), .Z(n138) );
  inv1f U77 ( .I(n87), .ZN(n66) );
  and2f U83 ( .A1(g0), .A2(n149), .Z(n148) );
  or2f U84 ( .A1(n150), .A2(n151), .Z(n149) );
  and2f U85 ( .A1(n152), .A2(n153), .Z(n151) );
  and2f U91 ( .A1(n309), .A2(o), .Z(n141) );
  and2f U114 ( .A1(t), .A2(n146), .Z(n87) );
  and2f U115 ( .A1(r), .A2(s), .Z(n146) );
  or2f U121 ( .A1(n173), .A2(n174), .Z(n92) );
  or2f U149 ( .A1(n206), .A2(n207), .Z(n205) );
  and2f U150 ( .A1(n208), .A2(n209), .Z(n207) );
  or2f U156 ( .A1(n130), .A2(n198), .Z(n196) );
  or2f U158 ( .A1(n215), .A2(n197), .Z(n218) );
  or2f U192 ( .A1(n246), .A2(n215), .Z(n198) );
  inv1f U193 ( .I(n247), .ZN(n215) );
  or2f U194 ( .A1(t), .A2(y), .Z(n247) );
  and2f U195 ( .A1(n305), .A2(n217), .Z(n246) );
  and2f U211 ( .A1(n254), .A2(n255), .Z(n253) );
  and2f U231 ( .A1(b), .A2(n277), .Z(n252) );
  buf0 U267 ( .I(n304), .Z(j0) );
  or2f U268 ( .A1(n142), .A2(n143), .Z(n137) );
  and2 U269 ( .A1(n130), .A2(m), .Z(n81) );
  and2 U270 ( .A1(n87), .A2(n144), .Z(n143) );
  inv1 U271 ( .I(n157), .ZN(n173) );
  or2 U272 ( .A1(n132), .A2(n133), .Z(n125) );
  and2f U273 ( .A1(n136), .A2(p), .Z(n134) );
  and2f U274 ( .A1(n92), .A2(n93), .Z(n71) );
  inv1 U275 ( .I(n104), .ZN(n91) );
  and2f U276 ( .A1(n155), .A2(n104), .Z(n154) );
  or2f U277 ( .A1(n95), .A2(n92), .Z(n104) );
  and2f U278 ( .A1(n91), .A2(g0), .Z(n82) );
  inv1 U279 ( .I(x), .ZN(n217) );
  inv1 U280 ( .I(r), .ZN(n130) );
  or2 U281 ( .A1(n201), .A2(n211), .Z(n222) );
  or2 U282 ( .A1(n125), .A2(n126), .Z(n124) );
  inv1 U283 ( .I(e), .ZN(n270) );
  and2 U284 ( .A1(n306), .A2(f), .Z(n272) );
  and2 U285 ( .A1(r), .A2(n), .Z(n69) );
  and2 U286 ( .A1(n275), .A2(n276), .Z(n264) );
  inv1 U287 ( .I(h), .ZN(n273) );
  or2 U288 ( .A1(n264), .A2(n265), .Z(n263) );
  or2 U289 ( .A1(n197), .A2(n198), .Z(n195) );
  or2 U290 ( .A1(c0), .A2(d0), .Z(n157) );
  inv1 U291 ( .I(t), .ZN(n140) );
  and2 U292 ( .A1(p), .A2(n166), .Z(n158) );
  or2 U293 ( .A1(q), .A2(n144), .Z(n112) );
  inv1 U294 ( .I(n84), .ZN(n83) );
  and2 U295 ( .A1(n61), .A2(n62), .Z(n60) );
  and2 U296 ( .A1(n70), .A2(n71), .Z(n61) );
  and2 U297 ( .A1(n63), .A2(n64), .Z(n62) );
  inv1 U298 ( .I(n112), .ZN(n86) );
  or2 U299 ( .A1(n281), .A2(n282), .Z(n280) );
  and2 U300 ( .A1(n291), .A2(n292), .Z(n289) );
  and2 U301 ( .A1(n216), .A2(n196), .Z(n212) );
  and2 U302 ( .A1(q), .A2(n171), .Z(n96) );
  or2 U303 ( .A1(n187), .A2(n188), .Z(n186) );
  and2 U304 ( .A1(p), .A2(n189), .Z(n188) );
  or2 U305 ( .A1(n252), .A2(n253), .Z(n250) );
  and2 U306 ( .A1(f0), .A2(n205), .Z(n204) );
  and2 U307 ( .A1(a), .A2(n147), .Z(n122) );
  or2 U308 ( .A1(n148), .A2(h0), .Z(n147) );
  and2 U309 ( .A1(n122), .A2(n123), .Z(r0) );
  or2f U310 ( .A1(n256), .A2(n257), .Z(n254) );
  or2 U311 ( .A1(h), .A2(n272), .Z(n271) );
  inv1 U312 ( .I(s), .ZN(n305) );
  inv1 U313 ( .I(s), .ZN(n131) );
  and2 U314 ( .A1(q), .A2(n131), .Z(n168) );
  inv1 U315 ( .I(d), .ZN(n306) );
  inv1 U316 ( .I(d), .ZN(n220) );
  or2 U317 ( .A1(e), .A2(n272), .Z(n274) );
  inv1 U318 ( .I(n272), .ZN(n265) );
  or2f U319 ( .A1(n293), .A2(n287), .Z(n291) );
  and2f U320 ( .A1(n280), .A2(n223), .Z(n279) );
  and2f U321 ( .A1(t), .A2(n163), .Z(n162) );
  or2f U322 ( .A1(n164), .A2(n165), .Z(n163) );
  or2f U323 ( .A1(n51), .A2(n50), .Z(n307) );
  and2f U324 ( .A1(n307), .A2(n308), .Z(s0) );
  and2 U325 ( .A1(a), .A2(n49), .Z(n308) );
  and2f U326 ( .A1(n87), .A2(n169), .Z(n161) );
  inv1f U327 ( .I(t), .ZN(n309) );
  and2 U328 ( .A1(n140), .A2(o), .Z(n310) );
  and2f U329 ( .A1(n138), .A2(n139), .Z(n311) );
  or2 U330 ( .A1(n140), .A2(n), .Z(n139) );
  and2f U331 ( .A1(n159), .A2(n160), .Z(n150) );
  or2f U332 ( .A1(n161), .A2(n162), .Z(n160) );
  and2f U333 ( .A1(n276), .A2(n220), .Z(n293) );
  and2f U334 ( .A1(d), .A2(n276), .Z(n286) );
  or2f U335 ( .A1(n270), .A2(n273), .Z(n276) );
  or2f U336 ( .A1(n170), .A2(n96), .Z(n169) );
  and2f U337 ( .A1(n69), .A2(p), .Z(n167) );
  and2f U338 ( .A1(n81), .A2(n158), .Z(n165) );
  inv1 U339 ( .I(n243), .ZN(n211) );
  and2 U340 ( .A1(n244), .A2(n200), .Z(n243) );
  or2 U341 ( .A1(p), .A2(u), .Z(n244) );
  inv1 U342 ( .I(i0), .ZN(n56) );
  inv1 U343 ( .I(h0), .ZN(n304) );
  inv1 U344 ( .I(c), .ZN(n223) );
  or2 U345 ( .A1(n217), .A2(n218), .Z(n216) );
  inv1 U346 ( .I(w), .ZN(n197) );
  or2 U347 ( .A1(n215), .A2(n131), .Z(n214) );
  and2 U348 ( .A1(q), .A2(n72), .Z(n70) );
  and2 U349 ( .A1(n71), .A2(n87), .Z(n85) );
  and2 U350 ( .A1(n94), .A2(n95), .Z(n93) );
  inv1 U351 ( .I(d0), .ZN(n226) );
  inv1 U352 ( .I(f0), .ZN(n95) );
  inv1 U353 ( .I(n219), .ZN(n183) );
  or2 U354 ( .A1(n223), .A2(n220), .Z(n236) );
  or2 U355 ( .A1(n298), .A2(n299), .Z(n297) );
  and2 U356 ( .A1(n301), .A2(n304), .Z(n298) );
  and2 U357 ( .A1(n300), .A2(n56), .Z(n299) );
  inv1 U358 ( .I(n301), .ZN(n300) );
  and2 U359 ( .A1(c), .A2(n220), .Z(n296) );
  or2 U360 ( .A1(d), .A2(n304), .Z(n302) );
  inv1 U361 ( .I(b), .ZN(n255) );
  inv1 U362 ( .I(c0), .ZN(n228) );
  and2 U363 ( .A1(d0), .A2(n228), .Z(n240) );
  and2 U364 ( .A1(c0), .A2(n226), .Z(n241) );
  and2 U365 ( .A1(n222), .A2(e0), .Z(n235) );
  and2 U366 ( .A1(n236), .A2(n237), .Z(n234) );
  or2 U367 ( .A1(n228), .A2(n226), .Z(n237) );
  and2 U368 ( .A1(n232), .A2(n233), .Z(n231) );
  and2 U369 ( .A1(c0), .A2(n174), .Z(n233) );
  and2 U370 ( .A1(n225), .A2(d0), .Z(n232) );
  and2 U371 ( .A1(n183), .A2(n95), .Z(n224) );
  and2 U372 ( .A1(n221), .A2(n222), .Z(n206) );
  and2 U373 ( .A1(n236), .A2(n222), .Z(n225) );
  and2 U374 ( .A1(z), .A2(n248), .Z(n184) );
  and2 U375 ( .A1(n49), .A2(b), .Z(n248) );
  and2 U376 ( .A1(n199), .A2(u), .Z(n187) );
  and2 U377 ( .A1(n192), .A2(n200), .Z(n199) );
  and2 U378 ( .A1(d), .A2(c), .Z(n185) );
  or2 U379 ( .A1(n179), .A2(n180), .Z(n178) );
  and2 U380 ( .A1(n181), .A2(n94), .Z(n180) );
  and2 U381 ( .A1(g0), .A2(n182), .Z(n179) );
  inv1 U382 ( .I(n181), .ZN(n182) );
  inv1 U383 ( .I(n184), .ZN(n177) );
  or2 U384 ( .A1(n127), .A2(n128), .Z(n126) );
  or2 U385 ( .A1(n304), .A2(n94), .Z(n127) );
  or2 U386 ( .A1(n115), .A2(n116), .Z(n98) );
  or2 U387 ( .A1(n120), .A2(n121), .Z(n115) );
  inv1 U388 ( .I(a0), .ZN(n49) );
  and2 U389 ( .A1(n88), .A2(n89), .Z(n52) );
  and2 U390 ( .A1(n96), .A2(n87), .Z(n88) );
  inv1 U391 ( .I(n275), .ZN(n287) );
  or2 U392 ( .A1(h), .A2(e), .Z(n275) );
  or2 U393 ( .A1(n286), .A2(n287), .Z(n284) );
  inv1 U394 ( .I(n276), .ZN(n283) );
  inv1 U395 ( .I(n81), .ZN(n113) );
  inv1 U396 ( .I(l), .ZN(n144) );
  inv1 U397 ( .I(q), .ZN(n78) );
  or2 U398 ( .A1(l), .A2(n66), .Z(n76) );
  or2 U399 ( .A1(t), .A2(o), .Z(n72) );
  and2 U400 ( .A1(n65), .A2(n66), .Z(n64) );
  and2 U401 ( .A1(n67), .A2(n68), .Z(n63) );
  or2 U402 ( .A1(r), .A2(m), .Z(n67) );
  or2 U403 ( .A1(s), .A2(n69), .Z(n68) );
  or2 U404 ( .A1(d), .A2(n275), .Z(n292) );
  and2 U405 ( .A1(n283), .A2(d), .Z(n290) );
  and2 U406 ( .A1(n283), .A2(n220), .Z(n282) );
  and2 U407 ( .A1(n284), .A2(n285), .Z(n281) );
  or2 U408 ( .A1(n220), .A2(n275), .Z(n285) );
  and2 U409 ( .A1(n223), .A2(g), .Z(n260) );
  and2 U410 ( .A1(n268), .A2(n269), .Z(n267) );
  or2 U411 ( .A1(n273), .A2(n274), .Z(n268) );
  or2 U412 ( .A1(n270), .A2(n271), .Z(n269) );
  and2 U413 ( .A1(n260), .A2(n263), .Z(n266) );
  or2 U414 ( .A1(n261), .A2(n262), .Z(n258) );
  and2 U415 ( .A1(n264), .A2(n265), .Z(n261) );
  inv1 U416 ( .I(n263), .ZN(n262) );
  or2 U417 ( .A1(n226), .A2(n227), .Z(n219) );
  or2 U418 ( .A1(n174), .A2(n228), .Z(n227) );
  or2 U419 ( .A1(n245), .A2(n198), .Z(n201) );
  and2 U420 ( .A1(n130), .A2(n197), .Z(n245) );
  and2 U421 ( .A1(n195), .A2(n196), .Z(n194) );
  and2 U422 ( .A1(q), .A2(s), .Z(n166) );
  and2 U423 ( .A1(p), .A2(n86), .Z(n170) );
  and2 U424 ( .A1(n167), .A2(n168), .Z(n164) );
  inv1 U425 ( .I(n80), .ZN(n114) );
  and2 U426 ( .A1(q), .A2(n113), .Z(n142) );
  or2 U427 ( .A1(n172), .A2(n91), .Z(n129) );
  and2 U428 ( .A1(n92), .A2(n95), .Z(n172) );
  or2 U429 ( .A1(n146), .A2(t), .Z(n65) );
  and2 U430 ( .A1(n113), .A2(n114), .Z(n111) );
  or2 U431 ( .A1(n78), .A2(n66), .Z(n108) );
  inv1 U432 ( .I(n145), .ZN(n102) );
  or2 U433 ( .A1(k), .A2(n108), .Z(n145) );
  inv1 U434 ( .I(p), .ZN(n110) );
  and2 U435 ( .A1(n223), .A2(d), .Z(n301) );
  or2 U436 ( .A1(n278), .A2(n279), .Z(n277) );
  and2 U437 ( .A1(c), .A2(n288), .Z(n278) );
  or2 U438 ( .A1(n289), .A2(n290), .Z(n288) );
  and2 U439 ( .A1(n258), .A2(n259), .Z(n257) );
  and2 U440 ( .A1(n266), .A2(n267), .Z(n256) );
  inv1 U441 ( .I(n260), .ZN(n259) );
  inv1 U442 ( .I(e0), .ZN(n174) );
  or2 U443 ( .A1(n210), .A2(n211), .Z(n209) );
  and2 U444 ( .A1(n212), .A2(n213), .Z(n210) );
  or2 U445 ( .A1(n197), .A2(n214), .Z(n213) );
  and2 U446 ( .A1(n219), .A2(n220), .Z(n208) );
  and2 U447 ( .A1(n219), .A2(n223), .Z(n221) );
  inv1 U448 ( .I(n201), .ZN(n192) );
  or2 U449 ( .A1(q), .A2(v), .Z(n200) );
  or2 U450 ( .A1(n190), .A2(n191), .Z(n189) );
  and2 U451 ( .A1(n192), .A2(q), .Z(n191) );
  and2 U452 ( .A1(v), .A2(n193), .Z(n190) );
  inv1 U453 ( .I(n194), .ZN(n193) );
  and2 U454 ( .A1(f0), .A2(n183), .Z(n181) );
  and2 U455 ( .A1(n154), .A2(r), .Z(n153) );
  or2 U456 ( .A1(f0), .A2(n156), .Z(n155) );
  and2 U457 ( .A1(n157), .A2(e0), .Z(n156) );
  and2 U458 ( .A1(n310), .A2(n158), .Z(n152) );
  inv1 U459 ( .I(n129), .ZN(n159) );
  inv1 U460 ( .I(g0), .ZN(n94) );
  or2 U461 ( .A1(n134), .A2(n135), .Z(n133) );
  and2 U462 ( .A1(n108), .A2(n110), .Z(n135) );
  and2 U463 ( .A1(n137), .A2(n114), .Z(n136) );
  or2 U464 ( .A1(n120), .A2(n102), .Z(n132) );
  or2 U465 ( .A1(n84), .A2(n129), .Z(n128) );
  and2 U466 ( .A1(n130), .A2(n131), .Z(n121) );
  inv1 U467 ( .I(n65), .ZN(n120) );
  and2 U468 ( .A1(n106), .A2(n107), .Z(n100) );
  or2 U469 ( .A1(p), .A2(n108), .Z(n107) );
  or2 U470 ( .A1(n109), .A2(n110), .Z(n106) );
  and2 U471 ( .A1(n111), .A2(n112), .Z(n109) );
  or2 U472 ( .A1(n102), .A2(n103), .Z(n101) );
  and2 U473 ( .A1(n104), .A2(n105), .Z(n103) );
  or2 U474 ( .A1(g0), .A2(f0), .Z(n105) );
  or2 U475 ( .A1(n117), .A2(n118), .Z(n116) );
  and2 U476 ( .A1(n119), .A2(n94), .Z(n117) );
  inv1 U477 ( .I(n92), .ZN(n119) );
  and2 U478 ( .A1(n110), .A2(k), .Z(n171) );
  and2 U479 ( .A1(n85), .A2(n86), .Z(n57) );
  and2 U480 ( .A1(n90), .A2(n56), .Z(n89) );
  or2 U481 ( .A1(n71), .A2(n82), .Z(n90) );
  or2 U482 ( .A1(n223), .A2(n302), .Z(n294) );
  or2 U483 ( .A1(n296), .A2(n297), .Z(n295) );
  and2 U484 ( .A1(n250), .A2(n251), .Z(n249) );
  inv1 U485 ( .I(j), .ZN(n251) );
  and2 U486 ( .A1(n184), .A2(n228), .Z(n242) );
  and2 U487 ( .A1(n184), .A2(n239), .Z(n238) );
  or2 U488 ( .A1(n240), .A2(n241), .Z(n239) );
  or2 U489 ( .A1(n230), .A2(n231), .Z(n229) );
  and2 U490 ( .A1(n234), .A2(n235), .Z(n230) );
  or2 U491 ( .A1(n203), .A2(n204), .Z(n202) );
  and2 U492 ( .A1(n224), .A2(n225), .Z(n203) );
  or2 U493 ( .A1(n177), .A2(n178), .Z(n176) );
  or2 U494 ( .A1(n185), .A2(n186), .Z(n175) );
  and2 U495 ( .A1(n124), .A2(n49), .Z(n123) );
  and2 U496 ( .A1(i0), .A2(n97), .Z(n50) );
  and2 U497 ( .A1(n294), .A2(n295), .Z(k0) );
  and2 U498 ( .A1(n249), .A2(i), .Z(l0) );
  and2 U499 ( .A1(n242), .A2(n225), .Z(m0) );
  and2 U500 ( .A1(n238), .A2(n225), .Z(n0) );
  and2 U501 ( .A1(n184), .A2(n229), .Z(o0) );
  and2 U502 ( .A1(n184), .A2(n202), .Z(p0) );
  or2 U503 ( .A1(n175), .A2(n176), .Z(q0) );
endmodule

