
module frg2 ( n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, 
        x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, 
        f3, e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, 
        n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, 
        v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, 
        d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, q0, p0, o0, n0, m0, l0, 
        k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, 
        q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, w9, v9, u9, t9, s9, 
        r9, q9, p9, o9, n9, m9, l9, k9, j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, 
        z8, y8, x8, w8, v8, u8, t8, s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, 
        h8, g8, f8, e8, d8, c8, b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, 
        p7, o7, n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, 
        x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, 
        f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, 
        n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, 
        v4, u4, t4, s4, r4, q4, p4, o4 );
  input n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3,
         v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3,
         e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2,
         n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1,
         w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1,
         f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, q0, p0, o0,
         n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v,
         u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9, j9, i9, h9, g9,
         f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8, s8, r8, q8, p8,
         o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8, b8, a8, z7, y7,
         x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, i7, h7,
         g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, q6,
         p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5,
         y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5,
         h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4,
         q4, p4, o4;
  wire   n1245, n39, n40, n62, n82, n102, n120, n121, n122, n123, n125, n126,
         n127, n218, n219, n221, n222, n223, n227, n229, n230, n234, n235,
         n236, n237, n238, n254, n255, n256, n257, n258, n259, n262, n263,
         n264, n286, n287, n288, n289, n290, n293, n294, n295, n334, n335,
         n336, n337, n338, n341, n342, n343, n375, n376, n377, n498, n568,
         n586, n632, n638, n639, n656, n657, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n694, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1025, n1026, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1036, n1037, n1038, n1039, n1041,
         n1042, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1063,
         n1064, n1065, n1066, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1246;

  and2 U22 ( .A1(n40), .A2(m0), .Z(z4) );
  and2 U47 ( .A1(n62), .A2(m0), .Z(y4) );
  and2 U72 ( .A1(n82), .A2(m0), .Z(x4) );
  and2 U96 ( .A1(n102), .A2(m0), .Z(w4) );
  and2 U115 ( .A1(n120), .A2(n694), .Z(v6) );
  and2 U116 ( .A1(n121), .A2(n122), .Z(n120) );
  or2 U117 ( .A1(n123), .A2(m1), .Z(n122) );
  and2 U118 ( .A1(p0), .A2(n1242), .Z(n123) );
  or2 U119 ( .A1(n125), .A2(n126), .Z(n121) );
  and2 U120 ( .A1(n127), .A2(m0), .Z(v4) );
  and2 U208 ( .A1(n218), .A2(n219), .Z(s4) );
  or2 U209 ( .A1(n696), .A2(n221), .Z(n219) );
  or2 U210 ( .A1(n222), .A2(n223), .Z(n221) );
  or2 U214 ( .A1(l0), .A2(a3), .Z(n227) );
  and2 U215 ( .A1(n229), .A2(n230), .Z(n222) );
  or2 U216 ( .A1(l0), .A2(i3), .Z(n230) );
  or2 U219 ( .A1(m0), .A2(q3), .Z(n218) );
  or2 U222 ( .A1(n235), .A2(n236), .Z(n234) );
  inv1 U223 ( .I(n237), .ZN(n236) );
  or2 U224 ( .A1(n238), .A2(n1), .Z(n237) );
  and2 U225 ( .A1(n1), .A2(n238), .Z(n235) );
  and2 U247 ( .A1(n255), .A2(n256), .Z(r4) );
  or2 U248 ( .A1(n696), .A2(n257), .Z(n256) );
  or2 U249 ( .A1(n258), .A2(n259), .Z(n257) );
  or2 U253 ( .A1(l0), .A2(b3), .Z(n262) );
  and2 U254 ( .A1(n263), .A2(n264), .Z(n258) );
  or2 U255 ( .A1(l0), .A2(j3), .Z(n264) );
  or2 U258 ( .A1(m0), .A2(r3), .Z(n255) );
  and2 U284 ( .A1(n286), .A2(n287), .Z(q4) );
  or2 U285 ( .A1(n696), .A2(n288), .Z(n287) );
  or2 U286 ( .A1(n289), .A2(n290), .Z(n288) );
  or2 U290 ( .A1(l0), .A2(c3), .Z(n293) );
  and2 U291 ( .A1(n294), .A2(n295), .Z(n289) );
  or2 U292 ( .A1(l0), .A2(k3), .Z(n295) );
  or2 U295 ( .A1(m0), .A2(s3), .Z(n286) );
  and2 U317 ( .A1(n694), .A2(n1244), .Z(p6) );
  and2 U332 ( .A1(n334), .A2(n335), .Z(p4) );
  or2 U333 ( .A1(n696), .A2(n336), .Z(n335) );
  or2 U334 ( .A1(n337), .A2(n338), .Z(n336) );
  or2 U338 ( .A1(l0), .A2(d3), .Z(n341) );
  and2 U339 ( .A1(n342), .A2(n343), .Z(n337) );
  or2 U340 ( .A1(l3), .A2(l0), .Z(n343) );
  or2 U344 ( .A1(m0), .A2(t3), .Z(n334) );
  and2 U383 ( .A1(n375), .A2(n376), .Z(n1245) );
  or2 U384 ( .A1(n377), .A2(i4), .Z(n376) );
  inv1 U385 ( .I(f1), .ZN(n377) );
  or2 U386 ( .A1(n238), .A2(f1), .Z(n375) );
  inv1 U387 ( .I(i4), .ZN(n238) );
  or2 U389 ( .A1(k4), .A2(n0), .Z(n254) );
  and2 U425 ( .A1(g1), .A2(n1221), .Z(l5) );
  and2 U446 ( .A1(t3), .A2(m0), .Z(k5) );
  and2 U474 ( .A1(s3), .A2(m0), .Z(j5) );
  and2 U493 ( .A1(m0), .A2(r3), .Z(i5) );
  and2 U514 ( .A1(m0), .A2(q3), .Z(h5) );
  and2 U535 ( .A1(p3), .A2(m0), .Z(g5) );
  and2 U568 ( .A1(o3), .A2(m0), .Z(f5) );
  and2 U587 ( .A1(n3), .A2(m0), .Z(e5) );
  and2 U605 ( .A1(m3), .A2(m0), .Z(d5) );
  inv1 U624 ( .I(l4), .ZN(n498) );
  and2 U625 ( .A1(n568), .A2(m0), .Z(c5) );
  and2 U651 ( .A1(n586), .A2(m0), .Z(b5) );
  or2 U746 ( .A1(k4), .A2(n126), .Z(n39) );
  inv1 U747 ( .I(m1), .ZN(n126) );
  and2 U749 ( .A1(n632), .A2(m0), .Z(a5) );
  and2 U759 ( .A1(n638), .A2(n781), .Z(u6) );
  inv1 U760 ( .I(n782), .ZN(n638) );
  and2 U761 ( .A1(n694), .A2(m1), .Z(n639) );
  buf0 U762 ( .I(n1222), .Z(o4) );
  buf0 U763 ( .I(u3), .Z(t4) );
  buf0 U764 ( .I(v3), .Z(u4) );
  buf0 U765 ( .I(m4), .Z(m5) );
  buf0 U766 ( .I(n1243), .Z(s5) );
  buf0 U767 ( .I(n1243), .Z(t5) );
  buf0 U768 ( .I(n1243), .Z(u5) );
  buf0 U769 ( .I(n1243), .Z(v5) );
  buf0 U770 ( .I(n1243), .Z(w5) );
  buf0 U771 ( .I(n1241), .Z(h6) );
  buf0 U772 ( .I(n1240), .Z(i6) );
  buf0 U773 ( .I(n1239), .Z(j6) );
  buf0 U774 ( .I(n1238), .Z(k6) );
  buf0 U775 ( .I(n1237), .Z(l6) );
  buf0 U776 ( .I(k4), .Z(m6) );
  buf0 U777 ( .I(n1245), .Z(n6) );
  buf0 U782 ( .I(n1121), .Z(n660) );
  or2 U783 ( .A1(n1121), .A2(n823), .Z(n661) );
  or2 U786 ( .A1(n1195), .A2(n1016), .Z(n662) );
  or2 U789 ( .A1(n785), .A2(n786), .Z(n665) );
  buf0 U790 ( .I(n1116), .Z(n666) );
  or2 U792 ( .A1(n1169), .A2(n1168), .Z(n668) );
  or2 U793 ( .A1(k1), .A2(l1), .Z(n669) );
  buf0 U795 ( .I(n1134), .Z(n671) );
  inv1 U798 ( .I(n673), .ZN(n1179) );
  inv1 U799 ( .I(n697), .ZN(n674) );
  or2 U801 ( .A1(n1195), .A2(n1022), .Z(n675) );
  or2 U803 ( .A1(n1246), .A2(n1195), .Z(n676) );
  inv1 U810 ( .I(n680), .ZN(n1007) );
  or2 U811 ( .A1(n679), .A2(n788), .Z(n681) );
  or2 U812 ( .A1(n679), .A2(n788), .Z(n682) );
  or2 U813 ( .A1(n1100), .A2(n788), .Z(n683) );
  or2 U814 ( .A1(n1100), .A2(n788), .Z(n684) );
  inv1 U818 ( .I(n691), .ZN(n689) );
  inv1 U819 ( .I(n691), .ZN(n690) );
  inv1 U821 ( .I(n1228), .ZN(n692) );
  inv1 U823 ( .I(n1228), .ZN(n694) );
  inv1 U825 ( .I(m0), .ZN(n696) );
  inv1 U826 ( .I(k0), .ZN(n732) );
  or2 U827 ( .A1(n732), .A2(l0), .Z(n905) );
  inv1 U828 ( .I(n905), .ZN(n907) );
  and2 U829 ( .A1(l0), .A2(n732), .Z(n697) );
  and2 U830 ( .A1(j3), .A2(n673), .Z(n699) );
  and2 U831 ( .A1(r3), .A2(n1179), .Z(n698) );
  or2 U832 ( .A1(n699), .A2(n698), .Z(n632) );
  and2 U833 ( .A1(k3), .A2(n673), .Z(n701) );
  and2 U834 ( .A1(s3), .A2(n1179), .Z(n700) );
  or2 U835 ( .A1(n701), .A2(n700), .Z(n586) );
  and2 U836 ( .A1(l3), .A2(n673), .Z(n703) );
  and2 U837 ( .A1(t3), .A2(n1179), .Z(n702) );
  or2 U838 ( .A1(n703), .A2(n702), .Z(n568) );
  and2 U839 ( .A1(d3), .A2(k0), .Z(n704) );
  or2 U840 ( .A1(n704), .A2(n907), .Z(n342) );
  and2 U841 ( .A1(n341), .A2(n732), .Z(n706) );
  inv1 U842 ( .I(l0), .ZN(n733) );
  or2 U843 ( .A1(n733), .A2(l3), .Z(n705) );
  and2 U844 ( .A1(n706), .A2(n705), .Z(n338) );
  inv1 U845 ( .I(o0), .ZN(n707) );
  inv1 U847 ( .I(b1), .ZN(n708) );
  and2 U848 ( .A1(l1), .A2(n708), .Z(n711) );
  inv1 U849 ( .I(a1), .ZN(n709) );
  and2 U850 ( .A1(k1), .A2(n709), .Z(n710) );
  or2 U851 ( .A1(n711), .A2(n710), .Z(n1158) );
  inv1 U852 ( .I(x0), .ZN(n712) );
  and2 U853 ( .A1(h1), .A2(n712), .Z(n715) );
  inv1 U854 ( .I(y0), .ZN(n713) );
  or2 U856 ( .A1(n715), .A2(n714), .Z(n718) );
  inv1 U857 ( .I(z0), .ZN(n716) );
  and2 U858 ( .A1(j1), .A2(n716), .Z(n717) );
  or2 U862 ( .A1(g4), .A2(h4), .Z(n720) );
  inv1 U863 ( .I(e4), .ZN(n1163) );
  and2 U867 ( .A1(n4), .A2(n1231), .Z(n721) );
  and2 U868 ( .A1(n1020), .A2(n721), .Z(n724) );
  and2 U870 ( .A1(d4), .A2(n1246), .Z(n722) );
  and2 U871 ( .A1(n1222), .A2(n722), .Z(n723) );
  or2 U872 ( .A1(n724), .A2(n723), .Z(n1244) );
  and2 U873 ( .A1(c3), .A2(k0), .Z(n725) );
  or2 U874 ( .A1(n725), .A2(n907), .Z(n294) );
  and2 U875 ( .A1(n293), .A2(n732), .Z(n727) );
  or2 U876 ( .A1(n733), .A2(k3), .Z(n726) );
  and2 U877 ( .A1(n727), .A2(n726), .Z(n290) );
  and2 U878 ( .A1(b3), .A2(k0), .Z(n728) );
  or2 U879 ( .A1(n728), .A2(n907), .Z(n263) );
  and2 U880 ( .A1(n262), .A2(n732), .Z(n730) );
  or2 U881 ( .A1(n733), .A2(j3), .Z(n729) );
  and2 U882 ( .A1(n730), .A2(n729), .Z(n259) );
  and2 U883 ( .A1(a3), .A2(k0), .Z(n731) );
  or2 U884 ( .A1(n731), .A2(n907), .Z(n229) );
  and2 U885 ( .A1(n227), .A2(n732), .Z(n735) );
  or2 U886 ( .A1(n733), .A2(i3), .Z(n734) );
  and2 U887 ( .A1(n735), .A2(n734), .Z(n223) );
  and2 U888 ( .A1(e3), .A2(n673), .Z(n737) );
  and2 U889 ( .A1(m3), .A2(n1179), .Z(n736) );
  or2 U890 ( .A1(n737), .A2(n736), .Z(n127) );
  inv1 U891 ( .I(n1244), .ZN(n125) );
  inv1 U892 ( .I(n0), .ZN(n1242) );
  and2 U893 ( .A1(f3), .A2(n673), .Z(n739) );
  and2 U894 ( .A1(n3), .A2(n1179), .Z(n738) );
  or2 U895 ( .A1(n739), .A2(n738), .Z(n102) );
  and2 U896 ( .A1(g3), .A2(n673), .Z(n741) );
  and2 U897 ( .A1(o3), .A2(n1179), .Z(n740) );
  or2 U898 ( .A1(n741), .A2(n740), .Z(n82) );
  and2 U899 ( .A1(h3), .A2(n673), .Z(n743) );
  and2 U900 ( .A1(p3), .A2(n1179), .Z(n742) );
  or2 U901 ( .A1(n743), .A2(n742), .Z(n62) );
  and2 U902 ( .A1(i3), .A2(n673), .Z(n745) );
  and2 U903 ( .A1(q3), .A2(n1179), .Z(n744) );
  or2 U904 ( .A1(n745), .A2(n744), .Z(n40) );
  inv1 U905 ( .I(h1), .ZN(n1241) );
  or2 U906 ( .A1(n1241), .A2(n254), .Z(n5) );
  inv1 U907 ( .I(i1), .ZN(n1240) );
  or2 U908 ( .A1(n1240), .A2(n254), .Z(o5) );
  inv1 U909 ( .I(j1), .ZN(n1239) );
  or2 U910 ( .A1(n1239), .A2(n254), .Z(p5) );
  or2 U912 ( .A1(n1238), .A2(n254), .Z(q5) );
  inv1 U913 ( .I(l1), .ZN(n1237) );
  or2 U914 ( .A1(n1237), .A2(n254), .Z(r5) );
  or2 U915 ( .A1(b4), .A2(c4), .Z(n748) );
  inv1 U916 ( .I(y3), .ZN(n1108) );
  or2 U918 ( .A1(n1108), .A2(n667), .Z(n746) );
  or2 U919 ( .A1(n746), .A2(a4), .Z(n747) );
  or2 U920 ( .A1(n748), .A2(n747), .Z(n749) );
  and2 U921 ( .A1(n749), .A2(n1), .Z(n751) );
  inv1 U922 ( .I(n749), .ZN(n1229) );
  and2 U923 ( .A1(n1245), .A2(n1229), .Z(n750) );
  or2 U924 ( .A1(n751), .A2(n750), .Z(n1243) );
  or2 U925 ( .A1(n1241), .A2(n39), .Z(x5) );
  or2 U926 ( .A1(n1240), .A2(n39), .Z(y5) );
  or2 U927 ( .A1(n1239), .A2(n39), .Z(z5) );
  or2 U928 ( .A1(n1238), .A2(n39), .Z(a6) );
  or2 U929 ( .A1(n1237), .A2(n39), .Z(b6) );
  or2 U930 ( .A1(n1241), .A2(n498), .Z(c6) );
  or2 U931 ( .A1(n1240), .A2(n498), .Z(d6) );
  or2 U932 ( .A1(n1239), .A2(n498), .Z(e6) );
  or2 U933 ( .A1(n1238), .A2(n498), .Z(f6) );
  or2 U934 ( .A1(n1237), .A2(n498), .Z(g6) );
  and2 U935 ( .A1(x3), .A2(n1229), .Z(o6) );
  or2 U936 ( .A1(d1), .A2(c1), .Z(n753) );
  or2 U941 ( .A1(n780), .A2(n1228), .Z(n752) );
  or2 U942 ( .A1(n753), .A2(n752), .Z(n754) );
  inv1 U943 ( .I(n754), .ZN(n757) );
  or2 U944 ( .A1(n1228), .A2(g1), .Z(n755) );
  inv1 U945 ( .I(n755), .ZN(n1194) );
  and2 U946 ( .A1(h1), .A2(n1194), .Z(n756) );
  or2 U947 ( .A1(n757), .A2(n756), .Z(q6) );
  or2 U948 ( .A1(c1), .A2(n671), .Z(n760) );
  and2 U949 ( .A1(g1), .A2(n780), .Z(n758) );
  or2 U950 ( .A1(n758), .A2(n1228), .Z(n766) );
  inv1 U951 ( .I(n766), .ZN(n759) );
  and2 U953 ( .A1(n1240), .A2(n780), .Z(n761) );
  inv1 U954 ( .I(n761), .ZN(n762) );
  inv1 U956 ( .I(d1), .ZN(n763) );
  or2 U957 ( .A1(n671), .A2(n763), .Z(n764) );
  and2 U958 ( .A1(n765), .A2(n764), .Z(r6) );
  or2 U959 ( .A1(n671), .A2(d1), .Z(n777) );
  and2 U960 ( .A1(n759), .A2(n777), .Z(n772) );
  and2 U961 ( .A1(n1239), .A2(n780), .Z(n767) );
  inv1 U962 ( .I(n767), .ZN(n770) );
  inv1 U963 ( .I(c1), .ZN(n768) );
  or2 U964 ( .A1(n671), .A2(n768), .Z(n769) );
  and2 U965 ( .A1(n770), .A2(n769), .Z(n771) );
  and2 U966 ( .A1(n772), .A2(n771), .Z(s6) );
  and2 U968 ( .A1(n1238), .A2(n780), .Z(n774) );
  inv1 U969 ( .I(n774), .ZN(n775) );
  and2 U970 ( .A1(n776), .A2(n775), .Z(t6) );
  or2 U971 ( .A1(n777), .A2(c1), .Z(n779) );
  or2 U972 ( .A1(g1), .A2(n1237), .Z(n778) );
  and2 U973 ( .A1(n779), .A2(n778), .Z(n782) );
  and2 U974 ( .A1(n694), .A2(n780), .Z(n781) );
  inv1 U980 ( .I(n665), .ZN(n1116) );
  inv1 U981 ( .I(n1134), .ZN(n788) );
  or2 U982 ( .A1(n679), .A2(n788), .Z(n898) );
  or2 U983 ( .A1(n681), .A2(n1), .Z(n787) );
  and2 U984 ( .A1(n694), .A2(n787), .Z(n792) );
  or2 U985 ( .A1(n1100), .A2(n788), .Z(n899) );
  or2 U986 ( .A1(n683), .A2(o1), .Z(n790) );
  or2 U987 ( .A1(n690), .A2(j0), .Z(n789) );
  and2 U988 ( .A1(n790), .A2(n789), .Z(n791) );
  and2 U989 ( .A1(n792), .A2(n791), .Z(w6) );
  or2 U990 ( .A1(n682), .A2(o1), .Z(n793) );
  and2 U991 ( .A1(n694), .A2(n793), .Z(n797) );
  or2 U992 ( .A1(n684), .A2(p1), .Z(n795) );
  or2 U993 ( .A1(n689), .A2(i0), .Z(n794) );
  and2 U994 ( .A1(n795), .A2(n794), .Z(n796) );
  and2 U995 ( .A1(n797), .A2(n796), .Z(x6) );
  or2 U996 ( .A1(n898), .A2(p1), .Z(n798) );
  and2 U997 ( .A1(n694), .A2(n798), .Z(n802) );
  or2 U998 ( .A1(n899), .A2(q1), .Z(n800) );
  or2 U999 ( .A1(n690), .A2(h0), .Z(n799) );
  and2 U1000 ( .A1(n800), .A2(n799), .Z(n801) );
  and2 U1001 ( .A1(n802), .A2(n801), .Z(y6) );
  or2 U1002 ( .A1(n681), .A2(q1), .Z(n803) );
  and2 U1003 ( .A1(n694), .A2(n803), .Z(n807) );
  or2 U1004 ( .A1(n683), .A2(r1), .Z(n805) );
  or2 U1005 ( .A1(n689), .A2(g0), .Z(n804) );
  and2 U1006 ( .A1(n805), .A2(n804), .Z(n806) );
  and2 U1007 ( .A1(n807), .A2(n806), .Z(z6) );
  or2 U1008 ( .A1(n682), .A2(r1), .Z(n808) );
  and2 U1009 ( .A1(n694), .A2(n808), .Z(n812) );
  or2 U1010 ( .A1(n684), .A2(s1), .Z(n810) );
  or2 U1011 ( .A1(n689), .A2(f0), .Z(n809) );
  and2 U1012 ( .A1(n810), .A2(n809), .Z(n811) );
  and2 U1013 ( .A1(n812), .A2(n811), .Z(a7) );
  or2 U1014 ( .A1(n898), .A2(s1), .Z(n813) );
  and2 U1015 ( .A1(n694), .A2(n813), .Z(n817) );
  or2 U1016 ( .A1(n899), .A2(t1), .Z(n815) );
  or2 U1017 ( .A1(n689), .A2(e0), .Z(n814) );
  and2 U1018 ( .A1(n815), .A2(n814), .Z(n816) );
  and2 U1019 ( .A1(n817), .A2(n816), .Z(b7) );
  or2 U1020 ( .A1(n681), .A2(t1), .Z(n818) );
  and2 U1021 ( .A1(n694), .A2(n818), .Z(n822) );
  or2 U1022 ( .A1(n683), .A2(u1), .Z(n820) );
  or2 U1023 ( .A1(n690), .A2(d0), .Z(n819) );
  and2 U1024 ( .A1(n820), .A2(n819), .Z(n821) );
  and2 U1025 ( .A1(n822), .A2(n821), .Z(c7) );
  or2 U1026 ( .A1(n0), .A2(m0), .Z(n823) );
  and2 U1027 ( .A1(n694), .A2(n1141), .Z(n827) );
  or2 U1028 ( .A1(n682), .A2(u1), .Z(n825) );
  or2 U1029 ( .A1(n684), .A2(v1), .Z(n824) );
  and2 U1030 ( .A1(n825), .A2(n824), .Z(n826) );
  and2 U1031 ( .A1(n827), .A2(n826), .Z(d7) );
  or2 U1032 ( .A1(n898), .A2(v1), .Z(n828) );
  and2 U1033 ( .A1(n694), .A2(n828), .Z(n832) );
  or2 U1034 ( .A1(n899), .A2(w1), .Z(n830) );
  or2 U1035 ( .A1(n690), .A2(k0), .Z(n829) );
  and2 U1036 ( .A1(n830), .A2(n829), .Z(n831) );
  and2 U1037 ( .A1(n832), .A2(n831), .Z(e7) );
  or2 U1038 ( .A1(n681), .A2(w1), .Z(n833) );
  and2 U1039 ( .A1(n694), .A2(n833), .Z(n837) );
  or2 U1040 ( .A1(n683), .A2(x1), .Z(n835) );
  or2 U1041 ( .A1(n689), .A2(l0), .Z(n834) );
  and2 U1042 ( .A1(n835), .A2(n834), .Z(n836) );
  and2 U1043 ( .A1(n837), .A2(n836), .Z(f7) );
  or2 U1044 ( .A1(n682), .A2(x1), .Z(n838) );
  and2 U1045 ( .A1(n694), .A2(n838), .Z(n842) );
  or2 U1046 ( .A1(n684), .A2(y1), .Z(n840) );
  or2 U1047 ( .A1(n689), .A2(q), .Z(n839) );
  and2 U1048 ( .A1(n840), .A2(n839), .Z(n841) );
  and2 U1049 ( .A1(n842), .A2(n841), .Z(g7) );
  or2 U1050 ( .A1(n898), .A2(y1), .Z(n843) );
  and2 U1051 ( .A1(n694), .A2(n843), .Z(n847) );
  or2 U1052 ( .A1(n899), .A2(z1), .Z(n845) );
  or2 U1053 ( .A1(n690), .A2(r), .Z(n844) );
  and2 U1054 ( .A1(n845), .A2(n844), .Z(n846) );
  and2 U1055 ( .A1(n847), .A2(n846), .Z(h7) );
  or2 U1056 ( .A1(n681), .A2(z1), .Z(n848) );
  and2 U1057 ( .A1(n694), .A2(n848), .Z(n852) );
  or2 U1058 ( .A1(n683), .A2(a2), .Z(n850) );
  or2 U1059 ( .A1(n689), .A2(s), .Z(n849) );
  and2 U1060 ( .A1(n850), .A2(n849), .Z(n851) );
  and2 U1061 ( .A1(n852), .A2(n851), .Z(i7) );
  or2 U1062 ( .A1(n682), .A2(a2), .Z(n853) );
  and2 U1063 ( .A1(n694), .A2(n853), .Z(n857) );
  or2 U1064 ( .A1(n684), .A2(b2), .Z(n855) );
  or2 U1065 ( .A1(n689), .A2(t), .Z(n854) );
  and2 U1066 ( .A1(n855), .A2(n854), .Z(n856) );
  and2 U1067 ( .A1(n857), .A2(n856), .Z(j7) );
  or2 U1068 ( .A1(n898), .A2(b2), .Z(n858) );
  and2 U1069 ( .A1(n694), .A2(n858), .Z(n862) );
  or2 U1070 ( .A1(n899), .A2(c2), .Z(n860) );
  or2 U1071 ( .A1(n689), .A2(u), .Z(n859) );
  and2 U1072 ( .A1(n860), .A2(n859), .Z(n861) );
  and2 U1073 ( .A1(n862), .A2(n861), .Z(k7) );
  or2 U1074 ( .A1(n681), .A2(c2), .Z(n863) );
  and2 U1075 ( .A1(n694), .A2(n863), .Z(n867) );
  or2 U1076 ( .A1(n683), .A2(d2), .Z(n865) );
  or2 U1077 ( .A1(n690), .A2(v), .Z(n864) );
  and2 U1078 ( .A1(n865), .A2(n864), .Z(n866) );
  and2 U1079 ( .A1(n867), .A2(n866), .Z(l7) );
  or2 U1080 ( .A1(n682), .A2(d2), .Z(n868) );
  and2 U1081 ( .A1(n694), .A2(n868), .Z(n872) );
  or2 U1082 ( .A1(n684), .A2(e2), .Z(n870) );
  or2 U1083 ( .A1(n689), .A2(w), .Z(n869) );
  and2 U1084 ( .A1(n870), .A2(n869), .Z(n871) );
  and2 U1085 ( .A1(n872), .A2(n871), .Z(m7) );
  or2 U1086 ( .A1(n898), .A2(e2), .Z(n873) );
  and2 U1087 ( .A1(n694), .A2(n873), .Z(n877) );
  or2 U1088 ( .A1(n899), .A2(f2), .Z(n875) );
  or2 U1089 ( .A1(n690), .A2(x), .Z(n874) );
  and2 U1090 ( .A1(n875), .A2(n874), .Z(n876) );
  and2 U1091 ( .A1(n877), .A2(n876), .Z(n7) );
  or2 U1092 ( .A1(n681), .A2(f2), .Z(n878) );
  and2 U1093 ( .A1(n692), .A2(n878), .Z(n882) );
  or2 U1094 ( .A1(n683), .A2(g2), .Z(n880) );
  or2 U1095 ( .A1(n690), .A2(y), .Z(n879) );
  and2 U1096 ( .A1(n880), .A2(n879), .Z(n881) );
  and2 U1097 ( .A1(n882), .A2(n881), .Z(o7) );
  or2 U1098 ( .A1(n682), .A2(g2), .Z(n883) );
  and2 U1099 ( .A1(n692), .A2(n883), .Z(n887) );
  or2 U1100 ( .A1(n684), .A2(h2), .Z(n885) );
  or2 U1101 ( .A1(n689), .A2(z), .Z(n884) );
  and2 U1102 ( .A1(n885), .A2(n884), .Z(n886) );
  and2 U1103 ( .A1(n887), .A2(n886), .Z(p7) );
  or2 U1104 ( .A1(n898), .A2(h2), .Z(n888) );
  and2 U1105 ( .A1(n692), .A2(n888), .Z(n892) );
  or2 U1106 ( .A1(n899), .A2(i2), .Z(n890) );
  or2 U1107 ( .A1(n690), .A2(a0), .Z(n889) );
  and2 U1108 ( .A1(n890), .A2(n889), .Z(n891) );
  and2 U1109 ( .A1(n892), .A2(n891), .Z(q7) );
  or2 U1110 ( .A1(n681), .A2(i2), .Z(n893) );
  and2 U1111 ( .A1(n692), .A2(n893), .Z(n897) );
  or2 U1112 ( .A1(n683), .A2(j2), .Z(n895) );
  or2 U1113 ( .A1(n689), .A2(b0), .Z(n894) );
  and2 U1114 ( .A1(n895), .A2(n894), .Z(n896) );
  and2 U1115 ( .A1(n897), .A2(n896), .Z(r7) );
  or2 U1116 ( .A1(n682), .A2(j2), .Z(n901) );
  or2 U1117 ( .A1(n684), .A2(k2), .Z(n900) );
  and2 U1118 ( .A1(n901), .A2(n900), .Z(n904) );
  or2 U1119 ( .A1(n690), .A2(c0), .Z(n902) );
  and2 U1120 ( .A1(n692), .A2(n902), .Z(n903) );
  and2 U1121 ( .A1(n904), .A2(n903), .Z(s7) );
  or2 U1123 ( .A1(n957), .A2(i), .Z(n906) );
  and2 U1124 ( .A1(n692), .A2(n906), .Z(n909) );
  or2 U1125 ( .A1(n1141), .A2(n907), .Z(n959) );
  or2 U1126 ( .A1(n959), .A2(a), .Z(n908) );
  and2 U1127 ( .A1(n909), .A2(n908), .Z(n914) );
  inv1 U1128 ( .I(n1141), .ZN(n910) );
  or2 U1129 ( .A1(n910), .A2(n1100), .Z(n962) );
  or2 U1130 ( .A1(n962), .A2(l2), .Z(n912) );
  or2 U1131 ( .A1(n910), .A2(n679), .Z(n963) );
  or2 U1132 ( .A1(n963), .A2(k2), .Z(n911) );
  and2 U1133 ( .A1(n912), .A2(n911), .Z(n913) );
  and2 U1134 ( .A1(n914), .A2(n913), .Z(t7) );
  or2 U1135 ( .A1(n957), .A2(j), .Z(n915) );
  and2 U1136 ( .A1(n692), .A2(n915), .Z(n917) );
  or2 U1137 ( .A1(n959), .A2(b), .Z(n916) );
  and2 U1138 ( .A1(n917), .A2(n916), .Z(n921) );
  or2 U1139 ( .A1(n962), .A2(m2), .Z(n919) );
  or2 U1140 ( .A1(n963), .A2(l2), .Z(n918) );
  and2 U1141 ( .A1(n919), .A2(n918), .Z(n920) );
  and2 U1142 ( .A1(n921), .A2(n920), .Z(u7) );
  or2 U1143 ( .A1(n957), .A2(k), .Z(n922) );
  and2 U1144 ( .A1(n692), .A2(n922), .Z(n924) );
  or2 U1145 ( .A1(n959), .A2(c), .Z(n923) );
  and2 U1146 ( .A1(n924), .A2(n923), .Z(n928) );
  or2 U1147 ( .A1(n962), .A2(n2), .Z(n926) );
  or2 U1148 ( .A1(n963), .A2(m2), .Z(n925) );
  and2 U1149 ( .A1(n926), .A2(n925), .Z(n927) );
  and2 U1150 ( .A1(n928), .A2(n927), .Z(v7) );
  or2 U1151 ( .A1(n957), .A2(l), .Z(n929) );
  and2 U1152 ( .A1(n692), .A2(n929), .Z(n931) );
  or2 U1153 ( .A1(n959), .A2(d), .Z(n930) );
  and2 U1154 ( .A1(n931), .A2(n930), .Z(n935) );
  or2 U1155 ( .A1(n962), .A2(o2), .Z(n933) );
  or2 U1156 ( .A1(n963), .A2(n2), .Z(n932) );
  and2 U1157 ( .A1(n933), .A2(n932), .Z(n934) );
  and2 U1158 ( .A1(n935), .A2(n934), .Z(w7) );
  or2 U1159 ( .A1(n957), .A2(m), .Z(n936) );
  and2 U1160 ( .A1(n692), .A2(n936), .Z(n938) );
  or2 U1161 ( .A1(n959), .A2(e), .Z(n937) );
  and2 U1162 ( .A1(n938), .A2(n937), .Z(n942) );
  or2 U1163 ( .A1(n962), .A2(p2), .Z(n940) );
  or2 U1164 ( .A1(n963), .A2(o2), .Z(n939) );
  and2 U1165 ( .A1(n940), .A2(n939), .Z(n941) );
  and2 U1166 ( .A1(n942), .A2(n941), .Z(x7) );
  or2 U1167 ( .A1(n957), .A2(n), .Z(n943) );
  and2 U1168 ( .A1(n692), .A2(n943), .Z(n945) );
  or2 U1169 ( .A1(n959), .A2(f), .Z(n944) );
  and2 U1170 ( .A1(n945), .A2(n944), .Z(n949) );
  or2 U1171 ( .A1(n962), .A2(q2), .Z(n947) );
  or2 U1172 ( .A1(n963), .A2(p2), .Z(n946) );
  and2 U1173 ( .A1(n947), .A2(n946), .Z(n948) );
  and2 U1174 ( .A1(n949), .A2(n948), .Z(y7) );
  or2 U1175 ( .A1(n957), .A2(o), .Z(n950) );
  and2 U1176 ( .A1(n692), .A2(n950), .Z(n952) );
  or2 U1177 ( .A1(n959), .A2(g), .Z(n951) );
  and2 U1178 ( .A1(n952), .A2(n951), .Z(n956) );
  or2 U1179 ( .A1(n962), .A2(r2), .Z(n954) );
  or2 U1180 ( .A1(n963), .A2(q2), .Z(n953) );
  and2 U1181 ( .A1(n954), .A2(n953), .Z(n955) );
  and2 U1182 ( .A1(n956), .A2(n955), .Z(z7) );
  or2 U1183 ( .A1(n957), .A2(p), .Z(n958) );
  and2 U1184 ( .A1(n692), .A2(n958), .Z(n961) );
  or2 U1185 ( .A1(n959), .A2(h), .Z(n960) );
  and2 U1186 ( .A1(n961), .A2(n960), .Z(n967) );
  or2 U1187 ( .A1(n962), .A2(s2), .Z(n965) );
  or2 U1188 ( .A1(n963), .A2(r2), .Z(n964) );
  and2 U1189 ( .A1(n965), .A2(n964), .Z(n966) );
  and2 U1190 ( .A1(n967), .A2(n966), .Z(a8) );
  or2 U1196 ( .A1(n971), .A2(n970), .Z(n973) );
  and2 U1197 ( .A1(n977), .A2(i), .Z(n972) );
  or2 U1198 ( .A1(n973), .A2(n972), .Z(n974) );
  and2 U1199 ( .A1(n694), .A2(n974), .Z(b8) );
  or2 U1202 ( .A1(n976), .A2(n975), .Z(n979) );
  inv1 U1203 ( .I(n1007), .ZN(n977) );
  and2 U1204 ( .A1(n977), .A2(j), .Z(n978) );
  or2 U1205 ( .A1(n979), .A2(n978), .Z(n980) );
  and2 U1206 ( .A1(n694), .A2(n980), .Z(c8) );
  or2 U1209 ( .A1(n982), .A2(n981), .Z(n984) );
  and2 U1210 ( .A1(n977), .A2(k), .Z(n983) );
  or2 U1211 ( .A1(n984), .A2(n983), .Z(n985) );
  and2 U1212 ( .A1(n694), .A2(n985), .Z(d8) );
  or2 U1215 ( .A1(n987), .A2(n986), .Z(n989) );
  and2 U1216 ( .A1(n977), .A2(l), .Z(n988) );
  or2 U1217 ( .A1(n989), .A2(n988), .Z(n990) );
  and2 U1218 ( .A1(n694), .A2(n990), .Z(e8) );
  or2 U1221 ( .A1(n992), .A2(n991), .Z(n994) );
  and2 U1222 ( .A1(n977), .A2(m), .Z(n993) );
  or2 U1223 ( .A1(n994), .A2(n993), .Z(n995) );
  and2 U1224 ( .A1(n694), .A2(n995), .Z(f8) );
  or2 U1227 ( .A1(n997), .A2(n996), .Z(n999) );
  and2 U1228 ( .A1(n977), .A2(n), .Z(n998) );
  or2 U1229 ( .A1(n999), .A2(n998), .Z(n1000) );
  and2 U1230 ( .A1(n694), .A2(n1000), .Z(g8) );
  or2 U1233 ( .A1(n1002), .A2(n1001), .Z(n1004) );
  and2 U1234 ( .A1(n977), .A2(o), .Z(n1003) );
  or2 U1235 ( .A1(n1004), .A2(n1003), .Z(n1005) );
  and2 U1236 ( .A1(n694), .A2(n1005), .Z(h8) );
  and2 U1237 ( .A1(z2), .A2(n1006), .Z(n1009) );
  and2 U1238 ( .A1(n977), .A2(p), .Z(n1008) );
  or2 U1239 ( .A1(n1009), .A2(n1008), .Z(n1010) );
  and2 U1240 ( .A1(n694), .A2(n1010), .Z(i8) );
  or2 U1241 ( .A1(n669), .A2(n1200), .Z(n1094) );
  inv1 U1242 ( .I(n1094), .ZN(n1011) );
  or2 U1243 ( .A1(n1011), .A2(n1241), .Z(n1021) );
  and2 U1244 ( .A1(l1), .A2(k1), .Z(n1015) );
  and2 U1245 ( .A1(j1), .A2(i1), .Z(n1013) );
  inv1 U1249 ( .I(k4), .ZN(n1155) );
  or2 U1250 ( .A1(n1155), .A2(n1246), .Z(n1016) );
  or2 U1251 ( .A1(n1020), .A2(n1016), .Z(n1198) );
  and2 U1254 ( .A1(a3), .A2(n686), .Z(n1026) );
  or2 U1255 ( .A1(n1155), .A2(n1228), .Z(n1019) );
  inv1 U1258 ( .I(n1021), .ZN(n1022) );
  and2 U1261 ( .A1(n1049), .A2(b3), .Z(n1025) );
  or2 U1262 ( .A1(n1026), .A2(n1025), .Z(j8) );
  and2 U1263 ( .A1(b3), .A2(n1097), .Z(n1029) );
  and2 U1265 ( .A1(n1046), .A2(c3), .Z(n1028) );
  or2 U1266 ( .A1(n1029), .A2(n1028), .Z(k8) );
  and2 U1267 ( .A1(c3), .A2(n685), .Z(n1032) );
  and2 U1269 ( .A1(n1030), .A2(d3), .Z(n1031) );
  or2 U1270 ( .A1(n1032), .A2(n1031), .Z(l8) );
  and2 U1271 ( .A1(d3), .A2(n1097), .Z(n1034) );
  and2 U1272 ( .A1(n1049), .A2(e3), .Z(n1033) );
  or2 U1273 ( .A1(n1034), .A2(n1033), .Z(m8) );
  and2 U1274 ( .A1(e3), .A2(n1097), .Z(n1037) );
  and2 U1276 ( .A1(n1030), .A2(f3), .Z(n1036) );
  or2 U1277 ( .A1(n1037), .A2(n1036), .Z(n8) );
  and2 U1278 ( .A1(f3), .A2(n1097), .Z(n1039) );
  and2 U1279 ( .A1(n1030), .A2(g3), .Z(n1038) );
  or2 U1280 ( .A1(n1039), .A2(n1038), .Z(o8) );
  and2 U1281 ( .A1(g3), .A2(n657), .Z(n1042) );
  and2 U1283 ( .A1(n1049), .A2(h3), .Z(n1041) );
  or2 U1284 ( .A1(n1042), .A2(n1041), .Z(p8) );
  and2 U1285 ( .A1(h3), .A2(n657), .Z(n1045) );
  and2 U1287 ( .A1(n1059), .A2(i3), .Z(n1044) );
  or2 U1288 ( .A1(n1045), .A2(n1044), .Z(q8) );
  and2 U1289 ( .A1(i3), .A2(n657), .Z(n1048) );
  or2 U1292 ( .A1(n1048), .A2(n1047), .Z(r8) );
  and2 U1293 ( .A1(j3), .A2(n685), .Z(n1051) );
  and2 U1295 ( .A1(n1049), .A2(k3), .Z(n1050) );
  or2 U1296 ( .A1(n1051), .A2(n1050), .Z(s8) );
  and2 U1297 ( .A1(k3), .A2(n685), .Z(n1054) );
  inv1 U1298 ( .I(n688), .ZN(n1052) );
  and2 U1299 ( .A1(n1052), .A2(l3), .Z(n1053) );
  or2 U1300 ( .A1(n1054), .A2(n1053), .Z(t8) );
  and2 U1301 ( .A1(l3), .A2(n686), .Z(n1056) );
  or2 U1303 ( .A1(n1056), .A2(n1055), .Z(u8) );
  and2 U1304 ( .A1(m3), .A2(n657), .Z(n1058) );
  and2 U1305 ( .A1(n1049), .A2(n3), .Z(n1057) );
  or2 U1306 ( .A1(n1058), .A2(n1057), .Z(v8) );
  and2 U1307 ( .A1(n3), .A2(n1097), .Z(n1061) );
  inv1 U1308 ( .I(n688), .ZN(n1059) );
  and2 U1309 ( .A1(n1059), .A2(o3), .Z(n1060) );
  or2 U1310 ( .A1(n1061), .A2(n1060), .Z(w8) );
  and2 U1311 ( .A1(o3), .A2(n685), .Z(n1064) );
  and2 U1313 ( .A1(n1030), .A2(p3), .Z(n1063) );
  or2 U1314 ( .A1(n1064), .A2(n1063), .Z(x8) );
  and2 U1315 ( .A1(p3), .A2(n657), .Z(n1066) );
  and2 U1316 ( .A1(n1049), .A2(q3), .Z(n1065) );
  or2 U1317 ( .A1(n1066), .A2(n1065), .Z(y8) );
  and2 U1318 ( .A1(q3), .A2(n685), .Z(n1069) );
  or2 U1321 ( .A1(n1069), .A2(n1068), .Z(z8) );
  and2 U1322 ( .A1(r3), .A2(n657), .Z(n1071) );
  and2 U1323 ( .A1(n1030), .A2(s3), .Z(n1070) );
  or2 U1324 ( .A1(n1071), .A2(n1070), .Z(a9) );
  and2 U1325 ( .A1(s3), .A2(n686), .Z(n1073) );
  and2 U1326 ( .A1(n1049), .A2(t3), .Z(n1072) );
  or2 U1327 ( .A1(n1073), .A2(n1072), .Z(b9) );
  and2 U1328 ( .A1(t3), .A2(n685), .Z(n1075) );
  or2 U1330 ( .A1(n1075), .A2(n1074), .Z(c9) );
  and2 U1331 ( .A1(u3), .A2(n685), .Z(n1077) );
  and2 U1332 ( .A1(n1030), .A2(v3), .Z(n1076) );
  or2 U1333 ( .A1(n1077), .A2(n1076), .Z(d9) );
  and2 U1334 ( .A1(v3), .A2(n1097), .Z(n1080) );
  and2 U1335 ( .A1(n1049), .A2(w3), .Z(n1079) );
  or2 U1336 ( .A1(n1080), .A2(n1079), .Z(e9) );
  inv1 U1337 ( .I(w0), .ZN(n1203) );
  or2 U1338 ( .A1(k1), .A2(n1203), .Z(n1081) );
  or2 U1339 ( .A1(n1081), .A2(n1200), .Z(n1091) );
  inv1 U1340 ( .I(t0), .ZN(n1082) );
  or2 U1341 ( .A1(j1), .A2(n1082), .Z(n1085) );
  inv1 U1342 ( .I(u0), .ZN(n1083) );
  or2 U1343 ( .A1(i1), .A2(n1083), .Z(n1084) );
  and2 U1344 ( .A1(n1085), .A2(n1084), .Z(n1086) );
  inv1 U1346 ( .I(v0), .ZN(n1199) );
  or2 U1347 ( .A1(n1200), .A2(n1199), .Z(n1087) );
  and2 U1348 ( .A1(n1088), .A2(n1087), .Z(n1089) );
  or2 U1349 ( .A1(n1089), .A2(l1), .Z(n1090) );
  inv1 U1352 ( .I(s0), .ZN(n1093) );
  or2 U1353 ( .A1(n1094), .A2(n1093), .Z(n1208) );
  and2 U1357 ( .A1(w3), .A2(n686), .Z(n1098) );
  or2 U1358 ( .A1(n1099), .A2(n1098), .Z(f9) );
  and2 U1359 ( .A1(x3), .A2(n1100), .Z(n1101) );
  or2 U1360 ( .A1(x3), .A2(n498), .Z(n1109) );
  or2 U1361 ( .A1(n1109), .A2(n666), .Z(n1104) );
  inv1 U1362 ( .I(n1104), .ZN(n1103) );
  or2 U1363 ( .A1(n1101), .A2(n1103), .Z(n1102) );
  and2 U1364 ( .A1(n689), .A2(n1102), .Z(g9) );
  or2 U1365 ( .A1(n1103), .A2(y3), .Z(n1106) );
  or2 U1366 ( .A1(n1104), .A2(n1108), .Z(n1105) );
  and2 U1367 ( .A1(n1106), .A2(n1105), .Z(n1107) );
  or2 U1368 ( .A1(n1107), .A2(n691), .Z(h9) );
  or2 U1369 ( .A1(n1109), .A2(n1108), .Z(n1117) );
  or2 U1370 ( .A1(n1117), .A2(n666), .Z(n1111) );
  inv1 U1371 ( .I(n1111), .ZN(n1110) );
  or2 U1372 ( .A1(n1110), .A2(z3), .Z(n1113) );
  or2 U1373 ( .A1(n1111), .A2(n667), .Z(n1112) );
  and2 U1374 ( .A1(n1113), .A2(n1112), .Z(n1114) );
  or2 U1375 ( .A1(n1114), .A2(n691), .Z(i9) );
  or2 U1376 ( .A1(n1116), .A2(n667), .Z(n1118) );
  and2 U1378 ( .A1(a4), .A2(n0), .Z(n1119) );
  and2 U1379 ( .A1(n1130), .A2(n1119), .Z(n1128) );
  and2 U1380 ( .A1(a4), .A2(n660), .Z(n1120) );
  inv1 U1382 ( .I(n660), .ZN(n1123) );
  and2 U1384 ( .A1(n1123), .A2(n1122), .Z(n1124) );
  or2 U1385 ( .A1(n1125), .A2(n1124), .Z(n1126) );
  inv1 U1390 ( .I(n1136), .ZN(n1131) );
  and2 U1391 ( .A1(n690), .A2(n1131), .Z(n1132) );
  or2 U1393 ( .A1(n671), .A2(n1228), .Z(n1180) );
  or2 U1394 ( .A1(n1180), .A2(n696), .Z(n1135) );
  inv1 U1395 ( .I(n1135), .ZN(n1191) );
  and2 U1396 ( .A1(b4), .A2(n1136), .Z(n1138) );
  inv1 U1398 ( .I(n1144), .ZN(n1137) );
  or2 U1401 ( .A1(n1191), .A2(n1140), .Z(k9) );
  or2 U1402 ( .A1(n1141), .A2(n1228), .Z(n1142) );
  inv1 U1403 ( .I(n1142), .ZN(n1182) );
  and2 U1405 ( .A1(n1144), .A2(n1143), .Z(n1145) );
  or2 U1406 ( .A1(n1182), .A2(n1145), .Z(l9) );
  and2 U1408 ( .A1(n1222), .A2(n1147), .Z(n1148) );
  or2 U1409 ( .A1(n1148), .A2(d4), .Z(n1152) );
  and2 U1410 ( .A1(n1194), .A2(n1198), .Z(n1150) );
  inv1 U1411 ( .I(d4), .ZN(n1149) );
  or2 U1412 ( .A1(n1150), .A2(n1149), .Z(n1151) );
  inv1 U1414 ( .I(n1180), .ZN(n1153) );
  or2 U1416 ( .A1(n691), .A2(g1), .Z(n1186) );
  or2 U1417 ( .A1(n1155), .A2(d4), .Z(n1156) );
  or2 U1418 ( .A1(n1246), .A2(n1156), .Z(n1162) );
  or2 U1419 ( .A1(n1159), .A2(n1158), .Z(n1160) );
  or2 U1421 ( .A1(n1162), .A2(n1161), .Z(n1164) );
  inv1 U1423 ( .I(n1164), .ZN(n1165) );
  or2 U1424 ( .A1(n1165), .A2(e4), .Z(n1166) );
  and2 U1425 ( .A1(n1169), .A2(n1166), .Z(n1167) );
  or2 U1426 ( .A1(n1186), .A2(n1167), .Z(n9) );
  or2 U1427 ( .A1(n664), .A2(n663), .Z(n1188) );
  inv1 U1428 ( .I(n1169), .ZN(n1170) );
  or2 U1429 ( .A1(n1170), .A2(f4), .Z(n1171) );
  and2 U1430 ( .A1(n668), .A2(n1171), .Z(n1172) );
  or2 U1431 ( .A1(n1172), .A2(n1186), .Z(o9) );
  inv1 U1432 ( .I(g4), .ZN(n1174) );
  inv1 U1434 ( .I(n1173), .ZN(n1177) );
  or2 U1437 ( .A1(n1177), .A2(n1176), .Z(n1178) );
  or2 U1439 ( .A1(n1180), .A2(n1179), .Z(n1181) );
  inv1 U1440 ( .I(n1181), .ZN(n1183) );
  or2 U1441 ( .A1(n1183), .A2(n1182), .Z(n1184) );
  or2 U1442 ( .A1(n1185), .A2(n1184), .Z(p9) );
  inv1 U1443 ( .I(n1186), .ZN(n1187) );
  and2 U1444 ( .A1(h4), .A2(n1187), .Z(n1190) );
  or2 U1445 ( .A1(n668), .A2(g4), .Z(n1189) );
  and2 U1446 ( .A1(n1190), .A2(n1189), .Z(n1192) );
  or2 U1447 ( .A1(n1192), .A2(n1191), .Z(q9) );
  and2 U1448 ( .A1(n234), .A2(n694), .Z(n1193) );
  and2 U1449 ( .A1(n679), .A2(n1193), .Z(r9) );
  and2 U1450 ( .A1(j4), .A2(n1194), .Z(n1220) );
  inv1 U1451 ( .I(n4), .ZN(n1196) );
  or2 U1452 ( .A1(n1196), .A2(n1195), .Z(n1197) );
  or2 U1453 ( .A1(n1198), .A2(n1197), .Z(n1218) );
  or2 U1454 ( .A1(n1199), .A2(n1238), .Z(n1202) );
  inv1 U1455 ( .I(n1200), .ZN(n1201) );
  and2 U1456 ( .A1(n1202), .A2(n1201), .Z(n1205) );
  or2 U1457 ( .A1(n1203), .A2(n1237), .Z(n1204) );
  and2 U1458 ( .A1(n1205), .A2(n1204), .Z(n1206) );
  or2 U1459 ( .A1(h1), .A2(n1206), .Z(n1207) );
  and2 U1460 ( .A1(n1208), .A2(n1207), .Z(n1216) );
  or2 U1461 ( .A1(h1), .A2(n669), .Z(n1210) );
  or2 U1462 ( .A1(u0), .A2(n1210), .Z(n1211) );
  and2 U1463 ( .A1(n1211), .A2(n1240), .Z(n1213) );
  and2 U1464 ( .A1(i1), .A2(t0), .Z(n1212) );
  or2 U1465 ( .A1(n1213), .A2(n1212), .Z(n1214) );
  inv1 U1466 ( .I(n1214), .ZN(n1215) );
  or2 U1467 ( .A1(n1216), .A2(n1215), .Z(n1217) );
  or2 U1468 ( .A1(n1218), .A2(n1217), .Z(n1219) );
  and2 U1469 ( .A1(n1220), .A2(n1219), .Z(n1227) );
  inv1 U1470 ( .I(j4), .ZN(n1221) );
  and2 U1471 ( .A1(n1221), .A2(n4), .Z(n1223) );
  inv1 U1472 ( .I(g1), .ZN(n1222) );
  and2 U1473 ( .A1(n1223), .A2(n1222), .Z(n1225) );
  and2 U1476 ( .A1(n1229), .A2(n639), .Z(t9) );
  and2 U1477 ( .A1(n1230), .A2(n639), .Z(u9) );
  and2 U1478 ( .A1(n1244), .A2(n694), .Z(n1234) );
  or2 U1479 ( .A1(n1232), .A2(n1231), .Z(n1233) );
  and2 U1480 ( .A1(n1234), .A2(n1233), .Z(v9) );
  inv1 U1481 ( .I(n1235), .ZN(w9) );
  inv1f U778 ( .I(n687), .ZN(n1049) );
  or2f U779 ( .A1(n673), .A2(m0), .Z(n1122) );
  or2f U780 ( .A1(n1133), .A2(n1132), .Z(j9) );
  inv1 U781 ( .I(n656), .ZN(n691) );
  and2 U784 ( .A1(n713), .A2(i1), .Z(n714) );
  inv1 U785 ( .I(f4), .ZN(n1168) );
  inv1 U787 ( .I(n1146), .ZN(n1147) );
  inv1 U788 ( .I(n1224), .ZN(n1099) );
  and2 U791 ( .A1(n1046), .A2(j3), .Z(n1047) );
  and2 U794 ( .A1(n1046), .A2(m3), .Z(n1055) );
  and2 U796 ( .A1(n1046), .A2(r3), .Z(n1068) );
  and2 U797 ( .A1(n1046), .A2(u3), .Z(n1074) );
  and2 U800 ( .A1(c4), .A2(n690), .Z(n1143) );
  or2f U802 ( .A1(n1128), .A2(n1127), .Z(n1129) );
  or2f U804 ( .A1(n1134), .A2(e1), .Z(n780) );
  and2f U805 ( .A1(n1018), .A2(n694), .Z(n686) );
  inv1 U806 ( .I(n1078), .ZN(n1030) );
  or2 U807 ( .A1(n1023), .A2(n1022), .Z(n688) );
  inv1 U808 ( .I(n1078), .ZN(n1046) );
  inv1f U809 ( .I(n969), .ZN(n678) );
  or2f U815 ( .A1(n1086), .A2(k1), .Z(n1088) );
  inv1f U816 ( .I(n968), .ZN(n1006) );
  and2f U817 ( .A1(n1018), .A2(n694), .Z(n657) );
  and2f U820 ( .A1(n1018), .A2(n694), .Z(n1097) );
  and2f U822 ( .A1(t2), .A2(n678), .Z(n970) );
  and2f U824 ( .A1(w2), .A2(n678), .Z(n986) );
  and2f U846 ( .A1(v2), .A2(n678), .Z(n981) );
  and2f U855 ( .A1(n760), .A2(n759), .Z(n773) );
  or2f U859 ( .A1(n1121), .A2(n0), .Z(n1134) );
  inv1f U860 ( .I(k1), .ZN(n1238) );
  inv1f U861 ( .I(n1231), .ZN(n1246) );
  and2f U864 ( .A1(x2), .A2(n678), .Z(n991) );
  and2f U865 ( .A1(y2), .A2(n678), .Z(n996) );
  and2f U866 ( .A1(u2), .A2(n678), .Z(n975) );
  and2f U869 ( .A1(z2), .A2(n678), .Z(n1001) );
  inv1f U911 ( .I(n1178), .ZN(n1185) );
  or2f U917 ( .A1(n668), .A2(n1174), .Z(n1173) );
  or2f U937 ( .A1(q0), .A2(n707), .Z(n1228) );
  and2f U938 ( .A1(v2), .A2(n1006), .Z(n987) );
  and2f U939 ( .A1(u2), .A2(n1006), .Z(n982) );
  and2f U940 ( .A1(x2), .A2(n1006), .Z(n997) );
  and2f U952 ( .A1(w2), .A2(n1006), .Z(n992) );
  and2f U955 ( .A1(n1200), .A2(n669), .Z(n1012) );
  or2f U967 ( .A1(i1), .A2(j1), .Z(n1200) );
  and2f U975 ( .A1(n1242), .A2(n1126), .Z(n1127) );
  or2f U976 ( .A1(n784), .A2(n1108), .Z(n785) );
  or2f U977 ( .A1(n1158), .A2(n1159), .Z(n1232) );
  or2f U978 ( .A1(n718), .A2(n717), .Z(n1159) );
  or2f U979 ( .A1(n1227), .A2(n1226), .Z(s9) );
  and2f U1122 ( .A1(n1091), .A2(n1090), .Z(n1092) );
  or2f U1191 ( .A1(k1), .A2(l1), .Z(n1209) );
  inv1f U1192 ( .I(n672), .ZN(n1141) );
  inv1f U1193 ( .I(n661), .ZN(n672) );
  or2f U1194 ( .A1(n905), .A2(n1141), .Z(n957) );
  or2f U1195 ( .A1(n1020), .A2(n1019), .Z(n1235) );
  inv1f U1200 ( .I(n1232), .ZN(n1020) );
  or2f U1201 ( .A1(a4), .A2(b4), .Z(n783) );
  and2f U1207 ( .A1(n690), .A2(n1139), .Z(n1140) );
  or2f U1208 ( .A1(n1138), .A2(n1137), .Z(n1139) );
  or2f U1213 ( .A1(n1136), .A2(b4), .Z(n1144) );
  or2 U1214 ( .A1(n1130), .A2(a4), .Z(n1136) );
  or2f U1219 ( .A1(n783), .A2(c4), .Z(n786) );
  or2f U1220 ( .A1(n1023), .A2(n1022), .Z(n1078) );
  and2f U1225 ( .A1(n773), .A2(n762), .Z(n765) );
  and2f U1226 ( .A1(n773), .A2(n777), .Z(n776) );
  and2f U1231 ( .A1(n1134), .A2(n692), .Z(n656) );
  or2f U1232 ( .A1(n1175), .A2(n1186), .Z(n1176) );
  and2f U1246 ( .A1(n1174), .A2(n1188), .Z(n1175) );
  or2f U1247 ( .A1(n1168), .A2(n1161), .Z(n664) );
  or2f U1248 ( .A1(n1161), .A2(n662), .Z(n1017) );
  and2f U1252 ( .A1(n672), .A2(n673), .Z(n680) );
  and2f U1253 ( .A1(y2), .A2(n1006), .Z(n1002) );
  and2f U1256 ( .A1(s2), .A2(n1006), .Z(n971) );
  and2f U1257 ( .A1(t2), .A2(n1006), .Z(n976) );
  and2f U1259 ( .A1(n905), .A2(n674), .Z(n673) );
  or2f U1260 ( .A1(n1235), .A2(n676), .Z(n1023) );
  inv1f U1264 ( .I(z3), .ZN(n667) );
  or2f U1268 ( .A1(n667), .A2(x3), .Z(n784) );
  inv1f U1275 ( .I(n679), .ZN(n1100) );
  and2f U1282 ( .A1(n1230), .A2(l4), .Z(n679) );
  or2f U1286 ( .A1(n785), .A2(n786), .Z(n1230) );
  and2f U1290 ( .A1(n1225), .A2(n1099), .Z(n1226) );
  and2f U1291 ( .A1(n1095), .A2(n1208), .Z(n1096) );
  or2f U1294 ( .A1(n1092), .A2(h1), .Z(n1095) );
  or2f U1302 ( .A1(n663), .A2(n1161), .Z(n1169) );
  inv1f U1312 ( .I(n1160), .ZN(n1161) );
  or2f U1319 ( .A1(n1162), .A2(n1163), .Z(n663) );
  or2f U1320 ( .A1(n720), .A2(n719), .Z(n1231) );
  or2f U1329 ( .A1(n1163), .A2(n1168), .Z(n719) );
  or2f U1345 ( .A1(n1154), .A2(n1153), .Z(m9) );
  and2f U1350 ( .A1(n1152), .A2(n1151), .Z(n1154) );
  or2f U1351 ( .A1(n1146), .A2(n675), .Z(n687) );
  or2f U1354 ( .A1(n1096), .A2(n1146), .Z(n1224) );
  or2f U1355 ( .A1(n1235), .A2(n1246), .Z(n1146) );
  or2f U1356 ( .A1(n1015), .A2(n1014), .Z(n1195) );
  or2f U1377 ( .A1(n1013), .A2(n1012), .Z(n1014) );
  and2f U1381 ( .A1(n1018), .A2(n694), .Z(n685) );
  or2f U1383 ( .A1(n1022), .A2(n1017), .Z(n1018) );
  and2f U1386 ( .A1(n694), .A2(n1129), .Z(n1133) );
  and2f U1387 ( .A1(n1130), .A2(n1120), .Z(n1125) );
  or2f U1388 ( .A1(n1118), .A2(n1117), .Z(n1130) );
  or2f U1389 ( .A1(n680), .A2(n1100), .Z(n969) );
  or2f U1392 ( .A1(n680), .A2(n679), .Z(n968) );
  or2f U1397 ( .A1(n677), .A2(n1200), .Z(n1121) );
  or2f U1399 ( .A1(n1209), .A2(h1), .Z(n677) );
endmodule

