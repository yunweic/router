
module i6 ( V133, V134, V97, V98, V99, V131, V96, V64, V32, V138, V205, V198, 
        V166 );
  input [1:0] V133;
  input [0:0] V134;
  input [0:0] V97;
  input [0:0] V98;
  input [0:0] V99;
  input [31:0] V131;
  input [31:0] V96;
  input [31:0] V64;
  input [31:0] V32;
  input [4:0] V138;
  output [6:0] V205;
  output [31:0] V198;
  output [27:0] V166;
  wire   V138_0, n1, n3, n251, n256, n261, n266, n271, n276, n281, n286, n291,
         n296, n301, n306, n311, n316, n321, n326, n331, n336, n341, n346,
         n351, n356, n361, n366, n371, n376, n381, n386, n389, n390, n391,
         n392, n393, n394, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n406, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n419, n420, n421, n423, n424, n425, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831;
  assign V138_0 = V138[0];

  and2 U1 ( .A1(V138[3]), .A2(n1), .Z(V205[6]) );
  and2 U3 ( .A1(V138_0), .A2(V134[0]), .Z(n3) );
  inv1 U286 ( .I(V64[9]), .ZN(n251) );
  inv1 U292 ( .I(V64[8]), .ZN(n256) );
  inv1 U298 ( .I(V64[7]), .ZN(n261) );
  inv1 U304 ( .I(V64[6]), .ZN(n266) );
  inv1 U310 ( .I(V64[5]), .ZN(n271) );
  inv1 U316 ( .I(V64[4]), .ZN(n276) );
  inv1 U322 ( .I(V64[3]), .ZN(n281) );
  inv1 U328 ( .I(V64[2]), .ZN(n286) );
  inv1 U334 ( .I(V64[27]), .ZN(n291) );
  inv1 U340 ( .I(V64[26]), .ZN(n296) );
  inv1 U346 ( .I(V64[25]), .ZN(n301) );
  inv1 U352 ( .I(V64[24]), .ZN(n306) );
  inv1 U358 ( .I(V64[23]), .ZN(n311) );
  inv1 U364 ( .I(V64[22]), .ZN(n316) );
  inv1 U370 ( .I(V64[21]), .ZN(n321) );
  inv1 U376 ( .I(V64[20]), .ZN(n326) );
  inv1 U382 ( .I(V64[1]), .ZN(n331) );
  inv1 U388 ( .I(V64[19]), .ZN(n336) );
  inv1 U394 ( .I(V64[18]), .ZN(n341) );
  inv1 U400 ( .I(V64[17]), .ZN(n346) );
  inv1 U406 ( .I(V64[16]), .ZN(n351) );
  inv1 U412 ( .I(V64[15]), .ZN(n356) );
  inv1 U418 ( .I(V64[14]), .ZN(n361) );
  inv1 U424 ( .I(V64[13]), .ZN(n366) );
  inv1 U430 ( .I(V64[12]), .ZN(n371) );
  inv1 U436 ( .I(V64[11]), .ZN(n376) );
  inv1 U442 ( .I(V64[10]), .ZN(n381) );
  inv1 U448 ( .I(V64[0]), .ZN(n386) );
  inv1 U457 ( .I(V138[2]), .ZN(n390) );
  inv1 U469 ( .I(V138[4]), .ZN(n401) );
  inv1 U477 ( .I(n394), .ZN(n409) );
  inv1 U478 ( .I(n394), .ZN(n410) );
  inv1 U483 ( .I(n542), .ZN(n415) );
  inv1 U484 ( .I(n542), .ZN(n416) );
  and2 U493 ( .A1(n413), .A2(V99[0]), .Z(n424) );
  or2 U494 ( .A1(n3), .A2(n424), .Z(n1) );
  and2 U495 ( .A1(n411), .A2(V32[0]), .Z(n430) );
  and2 U499 ( .A1(V64[0]), .A2(n410), .Z(n427) );
  or2 U500 ( .A1(n428), .A2(n427), .Z(n429) );
  or2 U501 ( .A1(n430), .A2(n429), .Z(V166[0]) );
  and2 U502 ( .A1(n826), .A2(V32[1]), .Z(n434) );
  and2 U504 ( .A1(V64[1]), .A2(n820), .Z(n431) );
  or2 U505 ( .A1(n432), .A2(n431), .Z(n433) );
  or2 U506 ( .A1(n434), .A2(n433), .Z(V166[1]) );
  and2 U507 ( .A1(n413), .A2(V32[2]), .Z(n438) );
  and2 U509 ( .A1(V64[2]), .A2(n820), .Z(n435) );
  or2 U510 ( .A1(n436), .A2(n435), .Z(n437) );
  or2 U511 ( .A1(n438), .A2(n437), .Z(V166[2]) );
  and2 U512 ( .A1(n412), .A2(V32[3]), .Z(n442) );
  and2 U513 ( .A1(n281), .A2(n818), .Z(n440) );
  and2 U514 ( .A1(V64[3]), .A2(n410), .Z(n439) );
  or2 U515 ( .A1(n440), .A2(n439), .Z(n441) );
  or2 U516 ( .A1(n442), .A2(n441), .Z(V166[3]) );
  and2 U517 ( .A1(n414), .A2(V32[4]), .Z(n446) );
  and2 U518 ( .A1(n276), .A2(n818), .Z(n444) );
  and2 U519 ( .A1(V64[4]), .A2(n409), .Z(n443) );
  or2 U521 ( .A1(n446), .A2(n445), .Z(V166[4]) );
  and2 U522 ( .A1(n411), .A2(V32[5]), .Z(n450) );
  and2 U523 ( .A1(n271), .A2(n817), .Z(n448) );
  and2 U524 ( .A1(V64[5]), .A2(n819), .Z(n447) );
  or2 U526 ( .A1(n450), .A2(n449), .Z(V166[5]) );
  and2 U527 ( .A1(n826), .A2(V32[6]), .Z(n454) );
  and2 U528 ( .A1(n266), .A2(n420), .Z(n452) );
  and2 U529 ( .A1(V64[6]), .A2(n820), .Z(n451) );
  or2 U531 ( .A1(n454), .A2(n453), .Z(V166[6]) );
  and2 U532 ( .A1(n413), .A2(V32[7]), .Z(n458) );
  and2 U533 ( .A1(n261), .A2(n420), .Z(n456) );
  and2 U534 ( .A1(V64[7]), .A2(n410), .Z(n455) );
  or2 U536 ( .A1(n458), .A2(n457), .Z(V166[7]) );
  and2 U537 ( .A1(n412), .A2(V32[8]), .Z(n462) );
  and2 U539 ( .A1(V64[8]), .A2(n409), .Z(n459) );
  or2 U540 ( .A1(n460), .A2(n459), .Z(n461) );
  or2 U541 ( .A1(n462), .A2(n461), .Z(V166[8]) );
  and2 U542 ( .A1(n414), .A2(V32[9]), .Z(n466) );
  and2 U544 ( .A1(V64[9]), .A2(n409), .Z(n463) );
  or2 U545 ( .A1(n464), .A2(n463), .Z(n465) );
  or2 U546 ( .A1(n466), .A2(n465), .Z(V166[9]) );
  and2 U547 ( .A1(n411), .A2(V32[10]), .Z(n470) );
  and2 U548 ( .A1(n381), .A2(n406), .Z(n468) );
  and2 U549 ( .A1(V64[10]), .A2(n819), .Z(n467) );
  or2 U551 ( .A1(n470), .A2(n469), .Z(V166[10]) );
  and2 U552 ( .A1(n826), .A2(V32[11]), .Z(n474) );
  and2 U553 ( .A1(n376), .A2(n421), .Z(n472) );
  and2 U554 ( .A1(V64[11]), .A2(n410), .Z(n471) );
  or2 U556 ( .A1(n474), .A2(n473), .Z(V166[11]) );
  and2 U557 ( .A1(n412), .A2(V32[12]), .Z(n478) );
  and2 U559 ( .A1(V64[12]), .A2(n819), .Z(n475) );
  or2 U560 ( .A1(n476), .A2(n475), .Z(n477) );
  or2 U561 ( .A1(n478), .A2(n477), .Z(V166[12]) );
  and2 U562 ( .A1(n414), .A2(V32[13]), .Z(n482) );
  and2 U563 ( .A1(n366), .A2(n406), .Z(n480) );
  and2 U564 ( .A1(V64[13]), .A2(n820), .Z(n479) );
  or2 U565 ( .A1(n480), .A2(n479), .Z(n481) );
  or2 U566 ( .A1(n482), .A2(n481), .Z(V166[13]) );
  and2 U567 ( .A1(n411), .A2(V32[14]), .Z(n486) );
  and2 U569 ( .A1(V64[14]), .A2(n409), .Z(n483) );
  or2 U570 ( .A1(n484), .A2(n483), .Z(n485) );
  or2 U571 ( .A1(n486), .A2(n485), .Z(V166[14]) );
  and2 U572 ( .A1(n826), .A2(V32[15]), .Z(n490) );
  and2 U574 ( .A1(V64[15]), .A2(n409), .Z(n487) );
  or2 U575 ( .A1(n488), .A2(n487), .Z(n489) );
  or2 U576 ( .A1(n490), .A2(n489), .Z(V166[15]) );
  and2 U577 ( .A1(n413), .A2(V32[16]), .Z(n494) );
  and2 U579 ( .A1(V64[16]), .A2(n409), .Z(n491) );
  or2 U580 ( .A1(n492), .A2(n491), .Z(n493) );
  or2 U581 ( .A1(n494), .A2(n493), .Z(V166[16]) );
  and2 U582 ( .A1(n412), .A2(V32[17]), .Z(n498) );
  and2 U584 ( .A1(V64[17]), .A2(n410), .Z(n495) );
  or2 U585 ( .A1(n496), .A2(n495), .Z(n497) );
  or2 U586 ( .A1(n498), .A2(n497), .Z(V166[17]) );
  and2 U587 ( .A1(n414), .A2(V32[18]), .Z(n502) );
  and2 U588 ( .A1(n341), .A2(n816), .Z(n500) );
  and2 U589 ( .A1(V64[18]), .A2(n409), .Z(n499) );
  or2 U590 ( .A1(n500), .A2(n499), .Z(n501) );
  or2 U591 ( .A1(n502), .A2(n501), .Z(V166[18]) );
  and2 U592 ( .A1(n411), .A2(V32[19]), .Z(n506) );
  and2 U593 ( .A1(n336), .A2(n823), .Z(n504) );
  and2 U594 ( .A1(V64[19]), .A2(n820), .Z(n503) );
  or2 U595 ( .A1(n504), .A2(n503), .Z(n505) );
  or2 U596 ( .A1(n506), .A2(n505), .Z(V166[19]) );
  and2 U597 ( .A1(n826), .A2(V32[20]), .Z(n510) );
  and2 U599 ( .A1(V64[20]), .A2(n820), .Z(n507) );
  or2 U600 ( .A1(n508), .A2(n507), .Z(n509) );
  or2 U601 ( .A1(n510), .A2(n509), .Z(V166[20]) );
  and2 U602 ( .A1(n413), .A2(V32[21]), .Z(n514) );
  and2 U604 ( .A1(V64[21]), .A2(n819), .Z(n511) );
  or2 U605 ( .A1(n512), .A2(n511), .Z(n513) );
  or2 U606 ( .A1(n514), .A2(n513), .Z(V166[21]) );
  and2 U607 ( .A1(n412), .A2(V32[22]), .Z(n518) );
  and2 U609 ( .A1(V64[22]), .A2(n820), .Z(n515) );
  or2 U610 ( .A1(n516), .A2(n515), .Z(n517) );
  or2 U611 ( .A1(n518), .A2(n517), .Z(V166[22]) );
  and2 U612 ( .A1(n414), .A2(V32[23]), .Z(n522) );
  and2 U614 ( .A1(V64[23]), .A2(n410), .Z(n519) );
  or2 U615 ( .A1(n520), .A2(n519), .Z(n521) );
  or2 U616 ( .A1(n522), .A2(n521), .Z(V166[23]) );
  and2 U617 ( .A1(n411), .A2(V32[24]), .Z(n526) );
  and2 U618 ( .A1(n306), .A2(n816), .Z(n524) );
  and2 U619 ( .A1(V64[24]), .A2(n410), .Z(n523) );
  or2 U620 ( .A1(n524), .A2(n523), .Z(n525) );
  or2 U621 ( .A1(n526), .A2(n525), .Z(V166[24]) );
  and2 U622 ( .A1(n826), .A2(V32[25]), .Z(n530) );
  and2 U624 ( .A1(V64[25]), .A2(n819), .Z(n527) );
  or2 U625 ( .A1(n528), .A2(n527), .Z(n529) );
  or2 U626 ( .A1(n530), .A2(n529), .Z(V166[25]) );
  and2 U627 ( .A1(n413), .A2(V32[26]), .Z(n534) );
  and2 U628 ( .A1(n296), .A2(n420), .Z(n532) );
  and2 U629 ( .A1(V64[26]), .A2(n819), .Z(n531) );
  or2 U631 ( .A1(n534), .A2(n533), .Z(V166[26]) );
  and2 U632 ( .A1(n412), .A2(V32[27]), .Z(n539) );
  and2 U633 ( .A1(n291), .A2(n420), .Z(n537) );
  and2 U634 ( .A1(V64[27]), .A2(n819), .Z(n536) );
  or2 U636 ( .A1(n539), .A2(n538), .Z(V166[27]) );
  and2 U637 ( .A1(V32[28]), .A2(V138[4]), .Z(n541) );
  and2 U638 ( .A1(n826), .A2(n541), .Z(n543) );
  or2 U639 ( .A1(n390), .A2(V138[4]), .Z(n542) );
  or2 U640 ( .A1(n543), .A2(n415), .Z(n548) );
  or2 U641 ( .A1(n421), .A2(V64[28]), .Z(n546) );
  inv1 U642 ( .I(V64[28]), .ZN(n544) );
  and2 U644 ( .A1(n546), .A2(n545), .Z(n547) );
  or2 U645 ( .A1(n548), .A2(n547), .Z(V198[0]) );
  and2 U646 ( .A1(V32[29]), .A2(V138[4]), .Z(n549) );
  and2 U647 ( .A1(n413), .A2(n549), .Z(n550) );
  or2 U648 ( .A1(n550), .A2(n822), .Z(n555) );
  inv1 U650 ( .I(V64[29]), .ZN(n551) );
  and2 U652 ( .A1(n553), .A2(n552), .Z(n554) );
  or2 U653 ( .A1(n555), .A2(n554), .Z(V198[1]) );
  and2 U654 ( .A1(V32[30]), .A2(V138[4]), .Z(n556) );
  and2 U655 ( .A1(n412), .A2(n556), .Z(n557) );
  or2 U656 ( .A1(n557), .A2(n415), .Z(n562) );
  or2 U657 ( .A1(n823), .A2(V64[30]), .Z(n560) );
  inv1 U658 ( .I(V64[30]), .ZN(n558) );
  and2 U660 ( .A1(n560), .A2(n559), .Z(n561) );
  or2 U661 ( .A1(n562), .A2(n561), .Z(V198[2]) );
  and2 U662 ( .A1(V32[31]), .A2(V138[4]), .Z(n563) );
  and2 U663 ( .A1(n414), .A2(n563), .Z(n564) );
  or2 U664 ( .A1(n564), .A2(n415), .Z(n569) );
  or2 U665 ( .A1(n828), .A2(V64[31]), .Z(n567) );
  inv1 U666 ( .I(V64[31]), .ZN(n565) );
  or2 U667 ( .A1(n417), .A2(n565), .Z(n566) );
  and2 U668 ( .A1(n567), .A2(n566), .Z(n568) );
  or2 U669 ( .A1(n569), .A2(n568), .Z(V198[3]) );
  and2 U670 ( .A1(V96[0]), .A2(V138[4]), .Z(n570) );
  and2 U671 ( .A1(n411), .A2(n570), .Z(n571) );
  or2 U672 ( .A1(n571), .A2(n415), .Z(n576) );
  or2 U673 ( .A1(n818), .A2(V131[0]), .Z(n574) );
  inv1 U674 ( .I(V131[0]), .ZN(n572) );
  or2 U675 ( .A1(n419), .A2(n572), .Z(n573) );
  and2 U676 ( .A1(n574), .A2(n573), .Z(n575) );
  or2 U677 ( .A1(n576), .A2(n575), .Z(V198[4]) );
  and2 U678 ( .A1(V96[1]), .A2(V138[4]), .Z(n577) );
  and2 U679 ( .A1(n826), .A2(n577), .Z(n578) );
  or2 U680 ( .A1(n578), .A2(n415), .Z(n583) );
  or2 U681 ( .A1(n816), .A2(V131[1]), .Z(n581) );
  inv1 U682 ( .I(V131[1]), .ZN(n579) );
  and2 U684 ( .A1(n581), .A2(n580), .Z(n582) );
  or2 U685 ( .A1(n583), .A2(n582), .Z(V198[5]) );
  and2 U686 ( .A1(V96[2]), .A2(V138[4]), .Z(n584) );
  and2 U687 ( .A1(n413), .A2(n584), .Z(n585) );
  or2 U688 ( .A1(n585), .A2(n415), .Z(n590) );
  or2 U689 ( .A1(n827), .A2(V131[2]), .Z(n588) );
  inv1 U690 ( .I(V131[2]), .ZN(n586) );
  or2 U691 ( .A1(n392), .A2(n586), .Z(n587) );
  and2 U692 ( .A1(n588), .A2(n587), .Z(n589) );
  and2 U694 ( .A1(V96[3]), .A2(V138[4]), .Z(n591) );
  and2 U695 ( .A1(n412), .A2(n591), .Z(n592) );
  or2 U696 ( .A1(n592), .A2(n416), .Z(n597) );
  or2 U697 ( .A1(n817), .A2(V131[3]), .Z(n595) );
  inv1 U698 ( .I(V131[3]), .ZN(n593) );
  or2 U699 ( .A1(n821), .A2(n593), .Z(n594) );
  and2 U700 ( .A1(n595), .A2(n594), .Z(n596) );
  or2 U701 ( .A1(n597), .A2(n596), .Z(V198[7]) );
  and2 U702 ( .A1(V96[4]), .A2(V138[4]), .Z(n598) );
  and2 U703 ( .A1(n414), .A2(n598), .Z(n599) );
  or2 U704 ( .A1(n599), .A2(n416), .Z(n604) );
  or2 U705 ( .A1(n421), .A2(V131[4]), .Z(n602) );
  inv1 U706 ( .I(V131[4]), .ZN(n600) );
  or2 U707 ( .A1(n417), .A2(n600), .Z(n601) );
  and2 U708 ( .A1(n602), .A2(n601), .Z(n603) );
  or2 U709 ( .A1(n604), .A2(n603), .Z(V198[8]) );
  and2 U710 ( .A1(V96[5]), .A2(V138[4]), .Z(n605) );
  and2 U711 ( .A1(n411), .A2(n605), .Z(n606) );
  or2 U712 ( .A1(n606), .A2(n415), .Z(n611) );
  or2 U713 ( .A1(n827), .A2(V131[5]), .Z(n609) );
  inv1 U714 ( .I(V131[5]), .ZN(n607) );
  or2 U715 ( .A1(n821), .A2(n607), .Z(n608) );
  and2 U716 ( .A1(n609), .A2(n608), .Z(n610) );
  or2 U717 ( .A1(n611), .A2(n610), .Z(V198[9]) );
  and2 U718 ( .A1(V96[6]), .A2(V138[4]), .Z(n612) );
  and2 U719 ( .A1(n414), .A2(n612), .Z(n613) );
  or2 U720 ( .A1(n613), .A2(n822), .Z(n618) );
  or2 U721 ( .A1(n828), .A2(V131[6]), .Z(n616) );
  inv1 U722 ( .I(V131[6]), .ZN(n614) );
  or2 U723 ( .A1(n419), .A2(n614), .Z(n615) );
  and2 U724 ( .A1(n616), .A2(n615), .Z(n617) );
  or2 U725 ( .A1(n618), .A2(n617), .Z(V198[10]) );
  and2 U726 ( .A1(V96[7]), .A2(V138[4]), .Z(n619) );
  and2 U727 ( .A1(n411), .A2(n619), .Z(n620) );
  or2 U728 ( .A1(n620), .A2(n415), .Z(n625) );
  or2 U729 ( .A1(n827), .A2(V131[7]), .Z(n623) );
  inv1 U730 ( .I(V131[7]), .ZN(n621) );
  or2 U731 ( .A1(n830), .A2(n621), .Z(n622) );
  and2 U732 ( .A1(n623), .A2(n622), .Z(n624) );
  or2 U733 ( .A1(n625), .A2(n624), .Z(V198[11]) );
  and2 U734 ( .A1(V96[8]), .A2(V138[4]), .Z(n626) );
  and2 U735 ( .A1(n412), .A2(n626), .Z(n627) );
  or2 U736 ( .A1(n627), .A2(n822), .Z(n632) );
  or2 U737 ( .A1(n420), .A2(V131[8]), .Z(n630) );
  inv1 U738 ( .I(V131[8]), .ZN(n628) );
  or2 U739 ( .A1(n392), .A2(n628), .Z(n629) );
  and2 U740 ( .A1(n630), .A2(n629), .Z(n631) );
  and2 U742 ( .A1(V96[9]), .A2(V138[4]), .Z(n633) );
  and2 U743 ( .A1(n826), .A2(n633), .Z(n634) );
  or2 U744 ( .A1(n634), .A2(n416), .Z(n639) );
  or2 U745 ( .A1(n818), .A2(V131[9]), .Z(n637) );
  inv1 U746 ( .I(V131[9]), .ZN(n635) );
  or2 U747 ( .A1(n821), .A2(n635), .Z(n636) );
  and2 U748 ( .A1(n637), .A2(n636), .Z(n638) );
  or2 U749 ( .A1(n638), .A2(n639), .Z(V198[13]) );
  and2 U750 ( .A1(V96[10]), .A2(V138[4]), .Z(n640) );
  and2 U751 ( .A1(n412), .A2(n640), .Z(n641) );
  or2 U752 ( .A1(n641), .A2(n415), .Z(n646) );
  or2 U753 ( .A1(n828), .A2(V131[10]), .Z(n644) );
  inv1 U754 ( .I(V131[10]), .ZN(n642) );
  and2 U756 ( .A1(n644), .A2(n643), .Z(n645) );
  or2 U757 ( .A1(n646), .A2(n645), .Z(V198[14]) );
  and2 U758 ( .A1(V96[11]), .A2(V138[4]), .Z(n647) );
  and2 U759 ( .A1(n414), .A2(n647), .Z(n648) );
  or2 U760 ( .A1(n648), .A2(n822), .Z(n653) );
  or2 U761 ( .A1(n816), .A2(V131[11]), .Z(n651) );
  inv1 U762 ( .I(V131[11]), .ZN(n649) );
  or2 U763 ( .A1(n392), .A2(n649), .Z(n650) );
  and2 U764 ( .A1(n651), .A2(n650), .Z(n652) );
  and2 U766 ( .A1(V96[12]), .A2(V138[4]), .Z(n654) );
  and2 U767 ( .A1(n826), .A2(n654), .Z(n655) );
  or2 U768 ( .A1(n655), .A2(n416), .Z(n660) );
  or2 U769 ( .A1(n421), .A2(V131[12]), .Z(n658) );
  inv1 U770 ( .I(V131[12]), .ZN(n656) );
  or2 U771 ( .A1(n830), .A2(n656), .Z(n657) );
  and2 U772 ( .A1(n658), .A2(n657), .Z(n659) );
  or2 U773 ( .A1(n660), .A2(n659), .Z(V198[16]) );
  and2 U774 ( .A1(V96[13]), .A2(V138[4]), .Z(n661) );
  and2 U775 ( .A1(n826), .A2(n661), .Z(n662) );
  or2 U776 ( .A1(n662), .A2(n822), .Z(n667) );
  or2 U777 ( .A1(n823), .A2(V131[13]), .Z(n665) );
  inv1 U778 ( .I(V131[13]), .ZN(n663) );
  and2 U780 ( .A1(n665), .A2(n664), .Z(n666) );
  or2 U781 ( .A1(n667), .A2(n666), .Z(V198[17]) );
  and2 U782 ( .A1(V96[14]), .A2(V138[4]), .Z(n668) );
  and2 U783 ( .A1(n413), .A2(n668), .Z(n669) );
  or2 U784 ( .A1(n669), .A2(n822), .Z(n674) );
  or2 U785 ( .A1(n827), .A2(V131[14]), .Z(n672) );
  inv1 U786 ( .I(V131[14]), .ZN(n670) );
  or2 U787 ( .A1(n830), .A2(n670), .Z(n671) );
  and2 U788 ( .A1(n672), .A2(n671), .Z(n673) );
  or2 U789 ( .A1(n674), .A2(n673), .Z(V198[18]) );
  and2 U790 ( .A1(V96[15]), .A2(V138[4]), .Z(n675) );
  and2 U791 ( .A1(n412), .A2(n675), .Z(n676) );
  or2 U792 ( .A1(n676), .A2(n416), .Z(n681) );
  or2 U793 ( .A1(n823), .A2(V131[15]), .Z(n679) );
  inv1 U794 ( .I(V131[15]), .ZN(n677) );
  or2 U795 ( .A1(n417), .A2(n677), .Z(n678) );
  and2 U796 ( .A1(n679), .A2(n678), .Z(n680) );
  or2 U797 ( .A1(n681), .A2(n680), .Z(V198[19]) );
  and2 U798 ( .A1(V96[16]), .A2(V138[4]), .Z(n682) );
  and2 U799 ( .A1(n412), .A2(n682), .Z(n683) );
  or2 U800 ( .A1(n683), .A2(n416), .Z(n688) );
  or2 U801 ( .A1(n406), .A2(V131[16]), .Z(n686) );
  inv1 U802 ( .I(V131[16]), .ZN(n684) );
  or2 U803 ( .A1(n419), .A2(n684), .Z(n685) );
  and2 U804 ( .A1(n686), .A2(n685), .Z(n687) );
  or2 U805 ( .A1(n688), .A2(n687), .Z(V198[20]) );
  and2 U806 ( .A1(V96[17]), .A2(V138[4]), .Z(n689) );
  and2 U807 ( .A1(n414), .A2(n689), .Z(n690) );
  or2 U808 ( .A1(n690), .A2(n416), .Z(n695) );
  or2 U809 ( .A1(n818), .A2(V131[17]), .Z(n693) );
  inv1 U810 ( .I(V131[17]), .ZN(n691) );
  or2 U811 ( .A1(n830), .A2(n691), .Z(n692) );
  and2 U812 ( .A1(n693), .A2(n692), .Z(n694) );
  or2 U813 ( .A1(n695), .A2(n694), .Z(V198[21]) );
  and2 U814 ( .A1(V96[18]), .A2(V138[4]), .Z(n696) );
  and2 U815 ( .A1(n412), .A2(n696), .Z(n697) );
  or2 U816 ( .A1(n697), .A2(n822), .Z(n702) );
  or2 U817 ( .A1(n421), .A2(V131[18]), .Z(n700) );
  inv1 U818 ( .I(V131[18]), .ZN(n698) );
  or2 U819 ( .A1(n821), .A2(n698), .Z(n699) );
  and2 U820 ( .A1(n700), .A2(n699), .Z(n701) );
  or2 U821 ( .A1(n702), .A2(n701), .Z(V198[22]) );
  and2 U822 ( .A1(V96[19]), .A2(V138[4]), .Z(n703) );
  and2 U823 ( .A1(n414), .A2(n703), .Z(n704) );
  or2 U824 ( .A1(n704), .A2(n822), .Z(n709) );
  or2 U825 ( .A1(n406), .A2(V131[19]), .Z(n707) );
  inv1 U826 ( .I(V131[19]), .ZN(n705) );
  or2 U827 ( .A1(n392), .A2(n705), .Z(n706) );
  and2 U828 ( .A1(n707), .A2(n706), .Z(n708) );
  and2 U830 ( .A1(V96[20]), .A2(V138[4]), .Z(n710) );
  and2 U831 ( .A1(n411), .A2(n710), .Z(n711) );
  or2 U832 ( .A1(n711), .A2(n416), .Z(n716) );
  or2 U833 ( .A1(n817), .A2(V131[20]), .Z(n714) );
  inv1 U834 ( .I(V131[20]), .ZN(n712) );
  or2 U835 ( .A1(n821), .A2(n712), .Z(n713) );
  and2 U836 ( .A1(n714), .A2(n713), .Z(n715) );
  or2 U837 ( .A1(n716), .A2(n715), .Z(V198[24]) );
  and2 U838 ( .A1(V96[21]), .A2(V138[4]), .Z(n717) );
  and2 U839 ( .A1(n411), .A2(n717), .Z(n718) );
  or2 U840 ( .A1(n718), .A2(n822), .Z(n723) );
  or2 U841 ( .A1(n818), .A2(V131[21]), .Z(n721) );
  inv1 U842 ( .I(V131[21]), .ZN(n719) );
  and2 U844 ( .A1(n721), .A2(n720), .Z(n722) );
  or2 U845 ( .A1(n723), .A2(n722), .Z(V198[25]) );
  and2 U846 ( .A1(V96[22]), .A2(V138[4]), .Z(n724) );
  and2 U847 ( .A1(n826), .A2(n724), .Z(n725) );
  or2 U848 ( .A1(n725), .A2(n415), .Z(n730) );
  or2 U849 ( .A1(n817), .A2(V131[22]), .Z(n728) );
  inv1 U850 ( .I(V131[22]), .ZN(n726) );
  or2 U851 ( .A1(n419), .A2(n726), .Z(n727) );
  and2 U852 ( .A1(n728), .A2(n727), .Z(n729) );
  or2 U853 ( .A1(n730), .A2(n729), .Z(V198[26]) );
  and2 U854 ( .A1(V96[23]), .A2(V138[4]), .Z(n731) );
  and2 U855 ( .A1(n412), .A2(n731), .Z(n732) );
  or2 U856 ( .A1(n732), .A2(n415), .Z(n737) );
  or2 U857 ( .A1(n817), .A2(V131[23]), .Z(n735) );
  inv1 U858 ( .I(V131[23]), .ZN(n733) );
  or2 U859 ( .A1(n417), .A2(n733), .Z(n734) );
  and2 U860 ( .A1(n735), .A2(n734), .Z(n736) );
  or2 U861 ( .A1(n737), .A2(n736), .Z(V198[27]) );
  and2 U862 ( .A1(V96[24]), .A2(V138[4]), .Z(n738) );
  and2 U863 ( .A1(n414), .A2(n738), .Z(n739) );
  or2 U864 ( .A1(n739), .A2(n416), .Z(n744) );
  or2 U865 ( .A1(n406), .A2(V131[24]), .Z(n742) );
  inv1 U866 ( .I(V131[24]), .ZN(n740) );
  and2 U868 ( .A1(n742), .A2(n741), .Z(n743) );
  or2 U869 ( .A1(n744), .A2(n743), .Z(V198[28]) );
  and2 U870 ( .A1(V96[25]), .A2(V138[4]), .Z(n745) );
  and2 U871 ( .A1(n411), .A2(n745), .Z(n746) );
  or2 U872 ( .A1(n746), .A2(n416), .Z(n751) );
  or2 U873 ( .A1(n406), .A2(V131[25]), .Z(n749) );
  inv1 U874 ( .I(V131[25]), .ZN(n747) );
  or2 U875 ( .A1(n417), .A2(n747), .Z(n748) );
  and2 U876 ( .A1(n749), .A2(n748), .Z(n750) );
  or2 U877 ( .A1(n751), .A2(n750), .Z(V198[29]) );
  and2 U878 ( .A1(V96[26]), .A2(V138[4]), .Z(n752) );
  and2 U879 ( .A1(n826), .A2(n752), .Z(n753) );
  or2 U880 ( .A1(n753), .A2(n822), .Z(n758) );
  or2 U881 ( .A1(n828), .A2(V131[26]), .Z(n756) );
  inv1 U882 ( .I(V131[26]), .ZN(n754) );
  or2 U883 ( .A1(n392), .A2(n754), .Z(n755) );
  and2 U884 ( .A1(n756), .A2(n755), .Z(n757) );
  and2 U886 ( .A1(V96[27]), .A2(V138[4]), .Z(n759) );
  and2 U887 ( .A1(n414), .A2(n759), .Z(n760) );
  or2 U888 ( .A1(n760), .A2(n822), .Z(n765) );
  or2 U889 ( .A1(n816), .A2(V131[27]), .Z(n763) );
  inv1 U890 ( .I(V131[27]), .ZN(n761) );
  and2 U892 ( .A1(n763), .A2(n762), .Z(n764) );
  or2 U893 ( .A1(n765), .A2(n764), .Z(V198[31]) );
  inv1 U894 ( .I(V131[28]), .ZN(n766) );
  or2 U895 ( .A1(n535), .A2(n766), .Z(n767) );
  or2 U897 ( .A1(n397), .A2(V131[28]), .Z(n768) );
  or2 U899 ( .A1(n390), .A2(V138[3]), .Z(n770) );
  inv1 U900 ( .I(n770), .ZN(n814) );
  or2 U901 ( .A1(n771), .A2(n814), .Z(n774) );
  and2 U902 ( .A1(V138[3]), .A2(V96[28]), .Z(n772) );
  and2 U903 ( .A1(n414), .A2(n772), .Z(n773) );
  or2 U904 ( .A1(n774), .A2(n773), .Z(V205[0]) );
  inv1 U905 ( .I(V131[29]), .ZN(n775) );
  or2 U906 ( .A1(n391), .A2(n775), .Z(n776) );
  and2 U907 ( .A1(V138[3]), .A2(n776), .Z(n778) );
  or2 U908 ( .A1(n816), .A2(V131[29]), .Z(n777) );
  and2 U911 ( .A1(V96[29]), .A2(V138[3]), .Z(n780) );
  and2 U912 ( .A1(n411), .A2(n780), .Z(n781) );
  or2 U913 ( .A1(n782), .A2(n781), .Z(V205[1]) );
  inv1 U914 ( .I(V131[30]), .ZN(n783) );
  or2 U915 ( .A1(n829), .A2(n783), .Z(n784) );
  and2 U916 ( .A1(V138[3]), .A2(n784), .Z(n786) );
  or2 U917 ( .A1(n406), .A2(V131[30]), .Z(n785) );
  and2 U920 ( .A1(V96[30]), .A2(V138[3]), .Z(n788) );
  and2 U921 ( .A1(n826), .A2(n788), .Z(n789) );
  or2 U922 ( .A1(n790), .A2(n789), .Z(V205[2]) );
  inv1 U923 ( .I(V131[31]), .ZN(n791) );
  or2 U924 ( .A1(n535), .A2(n791), .Z(n792) );
  and2 U925 ( .A1(V138[3]), .A2(n792), .Z(n794) );
  or2 U926 ( .A1(n816), .A2(V131[31]), .Z(n793) );
  and2 U929 ( .A1(V96[31]), .A2(V138[3]), .Z(n796) );
  and2 U930 ( .A1(n413), .A2(n796), .Z(n797) );
  or2 U931 ( .A1(n798), .A2(n797), .Z(V205[3]) );
  inv1 U932 ( .I(V133[0]), .ZN(n799) );
  or2 U933 ( .A1(n391), .A2(n799), .Z(n800) );
  and2 U934 ( .A1(V138[3]), .A2(n800), .Z(n802) );
  or2 U935 ( .A1(n823), .A2(V133[0]), .Z(n801) );
  and2 U938 ( .A1(V97[0]), .A2(V138[3]), .Z(n804) );
  and2 U939 ( .A1(n413), .A2(n804), .Z(n805) );
  or2 U940 ( .A1(n806), .A2(n805), .Z(V205[4]) );
  inv1 U941 ( .I(V133[1]), .ZN(n807) );
  or2 U942 ( .A1(n829), .A2(n807), .Z(n808) );
  and2 U943 ( .A1(V138[3]), .A2(n808), .Z(n810) );
  or2 U944 ( .A1(n818), .A2(V133[1]), .Z(n809) );
  and2 U946 ( .A1(V98[0]), .A2(V138[3]), .Z(n811) );
  and2 U947 ( .A1(n411), .A2(n811), .Z(n812) );
  or2 U949 ( .A1(n815), .A2(n814), .Z(V205[5]) );
  inv1f U456 ( .I(n425), .ZN(n823) );
  and2 U458 ( .A1(n286), .A2(n827), .Z(n436) );
  or2 U459 ( .A1(n444), .A2(n443), .Z(n445) );
  and2 U460 ( .A1(n251), .A2(n828), .Z(n464) );
  or2 U461 ( .A1(n468), .A2(n467), .Z(n469) );
  and2 U462 ( .A1(n361), .A2(n828), .Z(n484) );
  and2 U463 ( .A1(n326), .A2(n827), .Z(n508) );
  and2 U464 ( .A1(n316), .A2(n827), .Z(n516) );
  and2 U465 ( .A1(n311), .A2(n828), .Z(n520) );
  and2f U466 ( .A1(n346), .A2(n420), .Z(n496) );
  and2f U467 ( .A1(n356), .A2(n420), .Z(n488) );
  and2f U468 ( .A1(n321), .A2(n420), .Z(n512) );
  or2f U470 ( .A1(n420), .A2(V64[29]), .Z(n553) );
  inv1 U471 ( .I(V138_0), .ZN(n825) );
  or2f U472 ( .A1(n448), .A2(n447), .Z(n449) );
  or2f U473 ( .A1(n452), .A2(n451), .Z(n453) );
  or2f U474 ( .A1(n456), .A2(n455), .Z(n457) );
  or2f U475 ( .A1(n472), .A2(n471), .Z(n473) );
  and2f U476 ( .A1(n256), .A2(n817), .Z(n460) );
  and2f U479 ( .A1(n331), .A2(n817), .Z(n432) );
  and2f U480 ( .A1(n371), .A2(n817), .Z(n476) );
  and2f U481 ( .A1(n386), .A2(n421), .Z(n428) );
  and2f U482 ( .A1(n351), .A2(n421), .Z(n492) );
  and2f U485 ( .A1(n301), .A2(n421), .Z(n528) );
  or2f U486 ( .A1(n532), .A2(n531), .Z(n533) );
  or2f U487 ( .A1(n537), .A2(n536), .Z(n538) );
  or2f U488 ( .A1(n392), .A2(n558), .Z(n559) );
  or2f U489 ( .A1(n590), .A2(n589), .Z(V198[6]) );
  or2f U490 ( .A1(n632), .A2(n631), .Z(V198[12]) );
  or2f U491 ( .A1(n653), .A2(n652), .Z(V198[15]) );
  or2f U492 ( .A1(n709), .A2(n708), .Z(V198[23]) );
  or2f U496 ( .A1(n758), .A2(n757), .Z(V198[30]) );
  inv1 U497 ( .I(n824), .ZN(n831) );
  inv1 U498 ( .I(n403), .ZN(n396) );
  or2f U503 ( .A1(n831), .A2(n719), .Z(n720) );
  or2f U508 ( .A1(n831), .A2(n551), .Z(n552) );
  or2f U520 ( .A1(n831), .A2(n740), .Z(n741) );
  or2f U525 ( .A1(n831), .A2(n642), .Z(n643) );
  or2f U530 ( .A1(n396), .A2(n663), .Z(n664) );
  or2f U535 ( .A1(n396), .A2(n579), .Z(n580) );
  or2f U538 ( .A1(n396), .A2(n544), .Z(n545) );
  or2f U543 ( .A1(n396), .A2(n761), .Z(n762) );
  inv1f U550 ( .I(n423), .ZN(n420) );
  inv1f U555 ( .I(n425), .ZN(n816) );
  inv1f U558 ( .I(n824), .ZN(n830) );
  inv1f U568 ( .I(n423), .ZN(n817) );
  inv1f U573 ( .I(n403), .ZN(n419) );
  inv1f U578 ( .I(n425), .ZN(n818) );
  or2f U583 ( .A1(n400), .A2(V138[2]), .Z(n398) );
  inv1 U598 ( .I(n394), .ZN(n819) );
  inv1 U603 ( .I(n394), .ZN(n820) );
  inv1f U608 ( .I(n393), .ZN(n535) );
  inv1f U613 ( .I(n404), .ZN(n821) );
  inv1f U623 ( .I(n425), .ZN(n406) );
  inv1f U630 ( .I(n423), .ZN(n421) );
  inv1f U635 ( .I(n404), .ZN(n392) );
  inv1 U643 ( .I(n542), .ZN(n822) );
  or2f U649 ( .A1(n813), .A2(n812), .Z(n815) );
  and2f U651 ( .A1(n810), .A2(n809), .Z(n813) );
  or2f U659 ( .A1(n779), .A2(n814), .Z(n782) );
  and2f U683 ( .A1(n778), .A2(n777), .Z(n779) );
  or2f U693 ( .A1(n787), .A2(n814), .Z(n790) );
  and2f U741 ( .A1(n786), .A2(n785), .Z(n787) );
  or2f U755 ( .A1(n803), .A2(n814), .Z(n806) );
  and2f U765 ( .A1(n802), .A2(n801), .Z(n803) );
  inv1f U779 ( .I(n397), .ZN(n425) );
  and2f U829 ( .A1(n769), .A2(n768), .Z(n771) );
  and2f U843 ( .A1(V138[3]), .A2(n767), .Z(n769) );
  or2f U867 ( .A1(n399), .A2(V138[2]), .Z(n824) );
  or2f U885 ( .A1(n825), .A2(n401), .Z(n399) );
  or2f U891 ( .A1(n795), .A2(n814), .Z(n798) );
  and2f U896 ( .A1(n794), .A2(n793), .Z(n795) );
  inv1f U898 ( .I(V138_0), .ZN(n400) );
  inv1f U909 ( .I(n540), .ZN(n826) );
  inv1f U910 ( .I(n540), .ZN(n411) );
  inv1f U918 ( .I(n540), .ZN(n414) );
  inv1f U919 ( .I(n540), .ZN(n413) );
  inv1f U927 ( .I(n540), .ZN(n412) );
  or2f U928 ( .A1(V138[2]), .A2(V138_0), .Z(n540) );
  and2f U936 ( .A1(V138[2]), .A2(V138_0), .Z(n397) );
  inv1f U937 ( .I(n404), .ZN(n417) );
  or2f U945 ( .A1(n398), .A2(n401), .Z(n404) );
  inv1f U948 ( .I(n423), .ZN(n828) );
  inv1f U950 ( .I(n423), .ZN(n827) );
  inv1f U951 ( .I(n397), .ZN(n423) );
  or2f U952 ( .A1(V138[2]), .A2(n400), .Z(n394) );
  or2f U953 ( .A1(V138[2]), .A2(n402), .Z(n393) );
  inv1f U954 ( .I(V138_0), .ZN(n402) );
  and2f U955 ( .A1(n389), .A2(V138_0), .Z(n829) );
  and2f U956 ( .A1(n389), .A2(V138_0), .Z(n391) );
  inv1f U957 ( .I(V138[2]), .ZN(n389) );
  or2f U958 ( .A1(n399), .A2(V138[2]), .Z(n403) );
endmodule

