
module C5315_iscas ( v5, u5, t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, 
        h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, 
        p4, o4, n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, 
        x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, 
        f3, e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, 
        n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, 
        v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, 
        d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, 
        l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, 
        r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, o10, n10, m10, 
        l10, k10, j10, i10, h10, g10, f10, e10, d10, c10, b10, a10, z9, y9, x9, 
        w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9, j9, i9, h9, g9, f9, 
        e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8, s8, r8, q8, p8, o8, n8, 
        m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8, b8, a8, z7, y7, x7, w7, v7, 
        u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, 
        c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, 
        k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5 );
  input v5, u5, t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5,
         d5, c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4,
         m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3,
         v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3,
         e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2,
         n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1,
         w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1,
         f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0,
         o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x,
         w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output o10, n10, m10, l10, k10, j10, i10, h10, g10, f10, e10, d10, c10, b10,
         a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9,
         j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8,
         s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8,
         b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7,
         k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6,
         t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6,
         c6, b6, a6, z5, y5, x5, w5;
  wire   i5, v4, j3, i3, n1, l1, a, y7, s7, h7, v585, z585, n11, n12, n13, n14,
         n15, n16, n17, n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n105, n106,
         n109, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n169,
         n170, n171, n172, n173, n174, n175, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n321, n322, n324, n325, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n359, n360, n361, n362, n364, n365, n366,
         n368, n369, n373, n375, n376, n378, n380, n381, n382, n384, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n407, n408, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n441, n442, n443, n444, n446, n447,
         n448, n450, n451, n452, n453, n454, n455, n456, n457, n458, n469,
         n470, n471, n472, n473, n480, n481, n482, n483, n504, n507, n508,
         n509, n510, n512, n513, n514, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n588, n589,
         n590, n591, n592, n593, n594, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n629, n630, n631, n632, n644, n645, n646,
         n647, n648, n649, n651, n652, n653, n654, n655, n656, n657, n660,
         n661, n664, n665, n666, n667, n668, n669, n678, n691, n692, n725,
         n726, n727, n728, n729, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n775, n776, n777, n778, n779, n781, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n834, n835, n836, n837, n838, n839, n840, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n873, n879, n882, n883, n884, n885, n886,
         n887, n888, n889, n892, n893, n894, n895, n896, n898, n902, n903,
         n905, n909, n910, n911, n912, n927, n933, n934, n935, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1115, n1117,
         n1118, n1120, n1121, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1182, n1183, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1216, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1296, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1315, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1484, n1485, n1486, n1487, n1488, n1491, n1492, n1493,
         n1494, n1496, n1497, n1499, n1500, n1502, n1504, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1519, n1520, n1521, n1522,
         n1536, n1546, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, q7, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024;
  assign y5 = i5;
  assign u6 = v4;
  assign v6 = j3;
  assign d7 = j3;
  assign x5 = i3;
  assign w5 = n1;
  assign s6 = n1;
  assign r6 = l1;
  assign t6 = a;
  assign z6 = a;
  assign a7 = a;
  assign b7 = a;
  assign c7 = a;
  assign w7 = y7;
  assign p7 = s7;
  assign g7 = h7;
  assign z5 = v585;
  assign e6 = v585;
  assign f6 = v585;
  assign d6 = z585;
  assign w6 = z585;
  assign r7 = q7;

  or2 U1 ( .A1(n11), .A2(n12), .Z(z9) );
  or2 U2 ( .A1(n13), .A2(n14), .Z(n12) );
  and2 U3 ( .A1(n0), .A2(n15), .Z(n14) );
  and2 U4 ( .A1(m0), .A2(n16), .Z(n13) );
  or2 U5 ( .A1(n17), .A2(n18), .Z(n11) );
  and2 U6 ( .A1(n1987), .A2(n20), .Z(n18) );
  and2 U7 ( .A1(n1997), .A2(n22), .Z(n17) );
  or2 U8 ( .A1(n23), .A2(n24), .Z(z8) );
  or2 U9 ( .A1(n25), .A2(n26), .Z(n24) );
  and2 U10 ( .A1(y), .A2(n15), .Z(n26) );
  and2 U11 ( .A1(x), .A2(n16), .Z(n25) );
  or2 U12 ( .A1(n27), .A2(n28), .Z(n23) );
  and2 U13 ( .A1(n1987), .A2(n29), .Z(n28) );
  and2 U14 ( .A1(n1997), .A2(n30), .Z(n27) );
  inv1 U15 ( .I(n31), .ZN(z7) );
  inv1 U16 ( .I(v4), .ZN(z585) );
  or2 U17 ( .A1(n32), .A2(n33), .Z(y9) );
  or2 U18 ( .A1(n34), .A2(n35), .Z(n33) );
  and2 U19 ( .A1(r), .A2(n15), .Z(n35) );
  and2 U20 ( .A1(q), .A2(n16), .Z(n34) );
  or2 U21 ( .A1(n36), .A2(n37), .Z(n32) );
  and2 U22 ( .A1(n1987), .A2(n38), .Z(n37) );
  and2 U23 ( .A1(n1997), .A2(n39), .Z(n36) );
  or2 U24 ( .A1(n40), .A2(n41), .Z(y8) );
  or2 U25 ( .A1(n42), .A2(n43), .Z(n41) );
  and2 U26 ( .A1(e), .A2(n15), .Z(n43) );
  and2 U27 ( .A1(z), .A2(n16), .Z(n42) );
  or2 U28 ( .A1(n44), .A2(n45), .Z(n40) );
  and2 U29 ( .A1(n1987), .A2(n46), .Z(n45) );
  and2 U30 ( .A1(n1997), .A2(n47), .Z(n44) );
  or2 U31 ( .A1(n48), .A2(n49), .Z(x9) );
  or2 U32 ( .A1(n50), .A2(n51), .Z(n49) );
  and2 U33 ( .A1(o), .A2(n52), .Z(n51) );
  and2 U34 ( .A1(n53), .A2(n54), .Z(n50) );
  or2 U35 ( .A1(n55), .A2(n56), .Z(n48) );
  and2 U36 ( .A1(j0), .A2(n1981), .Z(n56) );
  and2 U37 ( .A1(n1982), .A2(n59), .Z(n55) );
  or2 U38 ( .A1(n60), .A2(n61), .Z(x8) );
  or2 U39 ( .A1(n62), .A2(n63), .Z(n61) );
  and2 U40 ( .A1(f), .A2(n15), .Z(n63) );
  and2 U41 ( .A1(a0), .A2(n16), .Z(n62) );
  or2 U42 ( .A1(n64), .A2(n65), .Z(n60) );
  and2 U43 ( .A1(n1987), .A2(n66), .Z(n65) );
  and2 U44 ( .A1(n1997), .A2(n67), .Z(n64) );
  or2 U45 ( .A1(n68), .A2(n69), .Z(x7) );
  or2 U46 ( .A1(y6), .A2(n70), .Z(x6) );
  inv1 U47 ( .I(m1), .ZN(n70) );
  or2 U48 ( .A1(n71), .A2(n72), .Z(w9) );
  or2 U49 ( .A1(n73), .A2(n74), .Z(n72) );
  and2 U50 ( .A1(n52), .A2(n0), .Z(n74) );
  and2 U51 ( .A1(n53), .A2(n20), .Z(n73) );
  or2 U52 ( .A1(n75), .A2(n76), .Z(n71) );
  and2 U53 ( .A1(n1981), .A2(m0), .Z(n76) );
  and2 U54 ( .A1(n1982), .A2(n22), .Z(n75) );
  or2 U55 ( .A1(n77), .A2(n78), .Z(w8) );
  or2 U56 ( .A1(n79), .A2(n80), .Z(n78) );
  and2 U57 ( .A1(n), .A2(n15), .Z(n80) );
  and2 U58 ( .A1(p), .A2(n16), .Z(n79) );
  or2 U59 ( .A1(n81), .A2(n82), .Z(n77) );
  and2 U60 ( .A1(n1987), .A2(n83), .Z(n82) );
  and2 U61 ( .A1(n1997), .A2(n84), .Z(n81) );
  or2 U65 ( .A1(n91), .A2(n92), .Z(v9) );
  or2 U66 ( .A1(n93), .A2(n94), .Z(n92) );
  and2 U67 ( .A1(n52), .A2(r), .Z(n94) );
  and2 U68 ( .A1(n53), .A2(n38), .Z(n93) );
  or2 U69 ( .A1(n95), .A2(n96), .Z(n91) );
  and2 U70 ( .A1(n1981), .A2(q), .Z(n96) );
  and2 U71 ( .A1(n1982), .A2(n39), .Z(n95) );
  or2 U72 ( .A1(n97), .A2(n98), .Z(v8) );
  or2 U73 ( .A1(n99), .A2(n100), .Z(n98) );
  and2 U74 ( .A1(n52), .A2(y), .Z(n100) );
  and2 U75 ( .A1(n53), .A2(n29), .Z(n99) );
  or2 U76 ( .A1(n101), .A2(n102), .Z(n97) );
  and2 U77 ( .A1(n1981), .A2(x), .Z(n102) );
  and2 U78 ( .A1(n1982), .A2(n30), .Z(n101) );
  or2 U80 ( .A1(n104), .A2(n105), .Z(n69) );
  and2 U81 ( .A1(n106), .A2(n1979), .Z(n104) );
  and2 U82 ( .A1(n2019), .A2(n109), .Z(n106) );
  inv1 U84 ( .I(u4), .ZN(v585) );
  or2 U85 ( .A1(n111), .A2(n112), .Z(u9) );
  or2 U86 ( .A1(n113), .A2(n114), .Z(n112) );
  and2 U87 ( .A1(o0), .A2(n52), .Z(n114) );
  and2 U88 ( .A1(n53), .A2(n115), .Z(n113) );
  or2 U89 ( .A1(n116), .A2(n117), .Z(n111) );
  and2 U90 ( .A1(p0), .A2(n1981), .Z(n117) );
  and2 U91 ( .A1(n1982), .A2(n118), .Z(n116) );
  or2 U92 ( .A1(n119), .A2(n120), .Z(u8) );
  or2 U93 ( .A1(n121), .A2(n122), .Z(n120) );
  and2 U94 ( .A1(n52), .A2(e), .Z(n122) );
  and2 U95 ( .A1(n53), .A2(n46), .Z(n121) );
  or2 U96 ( .A1(n123), .A2(n124), .Z(n119) );
  and2 U97 ( .A1(n1981), .A2(z), .Z(n124) );
  and2 U98 ( .A1(n1982), .A2(n47), .Z(n123) );
  or2 U99 ( .A1(n125), .A2(n126), .Z(t9) );
  or2 U100 ( .A1(n127), .A2(n128), .Z(n126) );
  and2 U101 ( .A1(o0), .A2(n15), .Z(n128) );
  and2 U102 ( .A1(p0), .A2(n16), .Z(n127) );
  or2 U103 ( .A1(n129), .A2(n130), .Z(n125) );
  and2 U104 ( .A1(n1987), .A2(n115), .Z(n130) );
  and2 U105 ( .A1(n1997), .A2(n118), .Z(n129) );
  or2 U106 ( .A1(n131), .A2(n132), .Z(t8) );
  or2 U107 ( .A1(n133), .A2(n134), .Z(n132) );
  and2 U108 ( .A1(f), .A2(n52), .Z(n134) );
  and2 U109 ( .A1(n53), .A2(n66), .Z(n133) );
  or2 U110 ( .A1(n135), .A2(n136), .Z(n131) );
  and2 U111 ( .A1(a0), .A2(n1981), .Z(n136) );
  and2 U112 ( .A1(n1982), .A2(n67), .Z(n135) );
  inv1 U113 ( .I(n54), .ZN(s9) );
  or2 U114 ( .A1(n137), .A2(n138), .Z(s8) );
  or2 U115 ( .A1(n139), .A2(n140), .Z(n138) );
  and2 U116 ( .A1(n), .A2(n52), .Z(n140) );
  and2 U117 ( .A1(n53), .A2(n83), .Z(n139) );
  or2 U118 ( .A1(n141), .A2(n142), .Z(n137) );
  and2 U119 ( .A1(p), .A2(n1981), .Z(n142) );
  and2 U120 ( .A1(n1982), .A2(n84), .Z(n141) );
  inv1 U121 ( .I(n20), .ZN(r9) );
  or2 U122 ( .A1(n143), .A2(n144), .Z(r8) );
  or2 U123 ( .A1(n145), .A2(n146), .Z(n144) );
  and2 U124 ( .A1(c2), .A2(n147), .Z(n146) );
  and2 U125 ( .A1(n148), .A2(n149), .Z(n145) );
  or2 U126 ( .A1(n150), .A2(n151), .Z(n143) );
  and2 U127 ( .A1(b2), .A2(n152), .Z(n151) );
  and2 U128 ( .A1(n153), .A2(n31), .Z(n150) );
  inv1 U129 ( .I(n38), .ZN(q9) );
  or2 U130 ( .A1(n154), .A2(n155), .Z(q8) );
  or2 U131 ( .A1(n156), .A2(n157), .Z(n155) );
  and2 U132 ( .A1(n158), .A2(c2), .Z(n157) );
  and2 U133 ( .A1(n159), .A2(n149), .Z(n156) );
  or2 U134 ( .A1(n160), .A2(n161), .Z(n154) );
  and2 U135 ( .A1(n162), .A2(b2), .Z(n161) );
  and2 U136 ( .A1(n163), .A2(n31), .Z(n160) );
  inv1 U140 ( .I(n169), .ZN(q6) );
  inv1 U141 ( .I(n115), .ZN(p9) );
  inv1 U142 ( .I(n170), .ZN(p8) );
  or2 U143 ( .A1(n171), .A2(n172), .Z(n170) );
  or2 U144 ( .A1(n173), .A2(n174), .Z(n172) );
  or2 U145 ( .A1(n175), .A2(n1998), .Z(n174) );
  or2 U146 ( .A1(n177), .A2(n178), .Z(n175) );
  or2 U147 ( .A1(n179), .A2(n180), .Z(n173) );
  or2 U148 ( .A1(n181), .A2(n182), .Z(n171) );
  or2 U149 ( .A1(n183), .A2(n184), .Z(n182) );
  or2 U150 ( .A1(n185), .A2(n186), .Z(n181) );
  and2 U151 ( .A1(n187), .A2(n188), .Z(s7) );
  and2 U152 ( .A1(n1979), .A2(n189), .Z(n188) );
  and2 U153 ( .A1(n190), .A2(n2019), .Z(n187) );
  or2 U154 ( .A1(h5), .A2(n191), .Z(p6) );
  inv1 U155 ( .I(k), .ZN(n191) );
  and2 U156 ( .A1(n192), .A2(n193), .Z(o9) );
  and2 U157 ( .A1(n194), .A2(n195), .Z(n193) );
  and2 U158 ( .A1(y4), .A2(n169), .Z(n195) );
  and2 U159 ( .A1(x4), .A2(f4), .Z(n169) );
  inv1 U160 ( .I(n196), .ZN(n194) );
  or2 U161 ( .A1(u7), .A2(j6), .Z(n196) );
  or2 U162 ( .A1(n197), .A2(n198), .Z(u7) );
  inv1 U163 ( .I(n199), .ZN(n198) );
  or2 U164 ( .A1(n200), .A2(n201), .Z(n199) );
  and2 U165 ( .A1(n201), .A2(n200), .Z(n197) );
  and2 U166 ( .A1(n202), .A2(n203), .Z(n200) );
  or2 U167 ( .A1(n204), .A2(l2), .Z(n203) );
  inv1 U168 ( .I(n205), .ZN(n204) );
  or2 U169 ( .A1(n205), .A2(n206), .Z(n202) );
  or2 U170 ( .A1(n207), .A2(n208), .Z(n205) );
  and2 U171 ( .A1(n209), .A2(n210), .Z(n208) );
  inv1 U172 ( .I(n211), .ZN(n210) );
  and2 U173 ( .A1(n211), .A2(n212), .Z(n207) );
  inv1 U174 ( .I(n209), .ZN(n212) );
  or2 U175 ( .A1(n213), .A2(n214), .Z(n209) );
  and2 U176 ( .A1(n215), .A2(n216), .Z(n214) );
  and2 U177 ( .A1(n217), .A2(a3), .Z(n213) );
  inv1 U178 ( .I(n215), .ZN(n217) );
  or2 U179 ( .A1(n218), .A2(n219), .Z(n215) );
  and2 U180 ( .A1(c3), .A2(n220), .Z(n219) );
  and2 U181 ( .A1(e3), .A2(n221), .Z(n218) );
  or2 U182 ( .A1(n222), .A2(n223), .Z(n211) );
  and2 U183 ( .A1(n224), .A2(n225), .Z(n223) );
  inv1 U184 ( .I(n226), .ZN(n225) );
  and2 U185 ( .A1(n226), .A2(n227), .Z(n222) );
  inv1 U186 ( .I(n224), .ZN(n227) );
  or2 U187 ( .A1(n228), .A2(n229), .Z(n224) );
  and2 U188 ( .A1(g3), .A2(n230), .Z(n229) );
  and2 U189 ( .A1(j2), .A2(n231), .Z(n228) );
  or2 U190 ( .A1(n232), .A2(n233), .Z(n226) );
  and2 U191 ( .A1(r2), .A2(n234), .Z(n233) );
  and2 U192 ( .A1(y2), .A2(n235), .Z(n232) );
  or2 U193 ( .A1(n236), .A2(n237), .Z(n201) );
  and2 U194 ( .A1(n2), .A2(n238), .Z(n237) );
  and2 U195 ( .A1(p2), .A2(n239), .Z(n236) );
  and2 U196 ( .A1(n240), .A2(n241), .Z(n192) );
  inv1 U197 ( .I(n242), .ZN(n241) );
  or2 U198 ( .A1(n8), .A2(t7), .Z(n242) );
  and2 U199 ( .A1(n243), .A2(n244), .Z(t7) );
  or2 U200 ( .A1(n245), .A2(n246), .Z(n244) );
  inv1 U201 ( .I(n247), .ZN(n243) );
  and2 U202 ( .A1(n246), .A2(n245), .Z(n247) );
  and2 U203 ( .A1(n248), .A2(n249), .Z(n245) );
  or2 U204 ( .A1(n250), .A2(k3), .Z(n249) );
  inv1 U205 ( .I(n251), .ZN(n250) );
  or2 U206 ( .A1(n251), .A2(n252), .Z(n248) );
  or2 U207 ( .A1(n253), .A2(n254), .Z(n251) );
  and2 U208 ( .A1(n255), .A2(n256), .Z(n254) );
  inv1 U209 ( .I(n257), .ZN(n256) );
  and2 U210 ( .A1(n257), .A2(n258), .Z(n253) );
  inv1 U211 ( .I(n255), .ZN(n258) );
  or2 U212 ( .A1(n259), .A2(n260), .Z(n255) );
  and2 U213 ( .A1(n261), .A2(n262), .Z(n260) );
  and2 U214 ( .A1(b4), .A2(n263), .Z(n259) );
  inv1 U215 ( .I(n261), .ZN(n263) );
  or2 U216 ( .A1(n264), .A2(n265), .Z(n261) );
  and2 U217 ( .A1(i3), .A2(n266), .Z(n265) );
  and2 U218 ( .A1(q3), .A2(n267), .Z(n264) );
  or2 U219 ( .A1(n268), .A2(n269), .Z(n257) );
  and2 U220 ( .A1(n270), .A2(n271), .Z(n269) );
  and2 U221 ( .A1(n272), .A2(v3), .Z(n268) );
  inv1 U222 ( .I(n270), .ZN(n272) );
  or2 U223 ( .A1(n273), .A2(n274), .Z(n270) );
  and2 U224 ( .A1(x3), .A2(n275), .Z(n274) );
  and2 U225 ( .A1(z3), .A2(n276), .Z(n273) );
  or2 U226 ( .A1(n277), .A2(n278), .Z(n246) );
  and2 U227 ( .A1(m3), .A2(n279), .Z(n278) );
  and2 U228 ( .A1(o3), .A2(n280), .Z(n277) );
  and2 U229 ( .A1(c6), .A2(n281), .Z(n240) );
  inv1 U230 ( .I(n282), .ZN(o8) );
  or2 U231 ( .A1(n283), .A2(n284), .Z(n282) );
  or2 U232 ( .A1(n285), .A2(n286), .Z(n284) );
  or2 U233 ( .A1(n287), .A2(n288), .Z(n286) );
  or2 U234 ( .A1(n289), .A2(n290), .Z(n287) );
  or2 U235 ( .A1(n291), .A2(n292), .Z(n285) );
  or2 U236 ( .A1(n293), .A2(n294), .Z(n283) );
  or2 U237 ( .A1(n295), .A2(n296), .Z(n294) );
  or2 U238 ( .A1(n297), .A2(n298), .Z(n293) );
  and2 U239 ( .A1(n299), .A2(n300), .Z(o7) );
  and2 U240 ( .A1(n301), .A2(n302), .Z(n300) );
  and2 U241 ( .A1(n303), .A2(n304), .Z(n302) );
  and2 U242 ( .A1(n305), .A2(n306), .Z(n303) );
  and2 U243 ( .A1(n307), .A2(n308), .Z(n301) );
  and2 U244 ( .A1(n309), .A2(n310), .Z(n299) );
  and2 U245 ( .A1(n311), .A2(n312), .Z(n310) );
  and2 U246 ( .A1(n313), .A2(n314), .Z(n309) );
  and2 U247 ( .A1(k1), .A2(n315), .Z(o6) );
  inv1 U248 ( .I(i5), .ZN(n315) );
  and2 U253 ( .A1(n2008), .A2(n324), .Z(n322) );
  and2 U254 ( .A1(d5), .A2(n325), .Z(n321) );
  inv1 U259 ( .I(n59), .ZN(n9) );
  and2 U260 ( .A1(n332), .A2(n333), .Z(n8) );
  or2 U261 ( .A1(n334), .A2(n335), .Z(n333) );
  inv1 U262 ( .I(n336), .ZN(n332) );
  and2 U263 ( .A1(n335), .A2(n334), .Z(n336) );
  and2 U264 ( .A1(n337), .A2(n338), .Z(n334) );
  inv1 U265 ( .I(n339), .ZN(n338) );
  and2 U266 ( .A1(n340), .A2(n341), .Z(n339) );
  or2 U267 ( .A1(n341), .A2(n340), .Z(n337) );
  or2 U268 ( .A1(n342), .A2(n343), .Z(n340) );
  and2 U269 ( .A1(n344), .A2(n345), .Z(n343) );
  inv1 U270 ( .I(n346), .ZN(n342) );
  or2 U271 ( .A1(n345), .A2(n344), .Z(n346) );
  or2 U272 ( .A1(n347), .A2(n348), .Z(n344) );
  and2 U273 ( .A1(n349), .A2(n350), .Z(n348) );
  inv1 U274 ( .I(n351), .ZN(n347) );
  or2 U275 ( .A1(n350), .A2(n349), .Z(n351) );
  and2 U280 ( .A1(n360), .A2(t3), .Z(n359) );
  and2 U281 ( .A1(n361), .A2(n362), .Z(n360) );
  or2 U282 ( .A1(n1980), .A2(n364), .Z(n362) );
  inv1 U283 ( .I(h3), .ZN(n364) );
  or2 U284 ( .A1(h3), .A2(n365), .Z(n361) );
  and2 U286 ( .A1(n368), .A2(n369), .Z(n366) );
  or2 U287 ( .A1(n1980), .A2(n231), .Z(n369) );
  inv1 U288 ( .I(g3), .ZN(n231) );
  or2 U289 ( .A1(g3), .A2(n365), .Z(n368) );
  or2 U294 ( .A1(n375), .A2(n376), .Z(n373) );
  and2 U295 ( .A1(n1996), .A2(n378), .Z(n376) );
  and2 U296 ( .A1(n1994), .A2(n380), .Z(n375) );
  or2 U297 ( .A1(n381), .A2(n382), .Z(n335) );
  and2 U298 ( .A1(n1993), .A2(n384), .Z(n382) );
  and2 U299 ( .A1(n1995), .A2(n386), .Z(n381) );
  and2 U300 ( .A1(n387), .A2(n388), .Z(n7) );
  and2 U301 ( .A1(n389), .A2(n390), .Z(n388) );
  and2 U302 ( .A1(n391), .A2(n392), .Z(n390) );
  and2 U303 ( .A1(n393), .A2(n394), .Z(n391) );
  and2 U304 ( .A1(n395), .A2(n396), .Z(n389) );
  and2 U305 ( .A1(n397), .A2(n398), .Z(n387) );
  and2 U306 ( .A1(n399), .A2(n400), .Z(n398) );
  and2 U307 ( .A1(n401), .A2(n402), .Z(n397) );
  and2 U308 ( .A1(d4), .A2(a), .Z(n6) );
  and2 U313 ( .A1(n2010), .A2(n324), .Z(n408) );
  inv1 U314 ( .I(z1), .ZN(n324) );
  and2 U315 ( .A1(b5), .A2(n325), .Z(n407) );
  inv1 U316 ( .I(a2), .ZN(n325) );
  inv1 U324 ( .I(n22), .ZN(m9) );
  inv1 U325 ( .I(n281), .ZN(m8) );
  or2 U326 ( .A1(n416), .A2(n417), .Z(n281) );
  inv1 U327 ( .I(n418), .ZN(n417) );
  or2 U328 ( .A1(n419), .A2(n420), .Z(n418) );
  and2 U329 ( .A1(n420), .A2(n419), .Z(n416) );
  and2 U330 ( .A1(n421), .A2(n422), .Z(n419) );
  or2 U331 ( .A1(n423), .A2(n1984), .Z(n422) );
  inv1 U332 ( .I(n424), .ZN(n423) );
  or2 U333 ( .A1(n424), .A2(n425), .Z(n421) );
  or2 U334 ( .A1(n426), .A2(n427), .Z(n424) );
  and2 U335 ( .A1(n428), .A2(n429), .Z(n427) );
  inv1 U336 ( .I(n430), .ZN(n426) );
  or2 U337 ( .A1(n429), .A2(n428), .Z(n430) );
  or2 U338 ( .A1(n431), .A2(n432), .Z(n428) );
  and2 U339 ( .A1(n433), .A2(n434), .Z(n432) );
  inv1 U340 ( .I(n435), .ZN(n431) );
  or2 U341 ( .A1(n434), .A2(n433), .Z(n435) );
  and2 U346 ( .A1(n442), .A2(s3), .Z(n441) );
  and2 U347 ( .A1(n443), .A2(n444), .Z(n442) );
  or2 U348 ( .A1(n1999), .A2(n446), .Z(n444) );
  inv1 U349 ( .I(c4), .ZN(n446) );
  or2 U350 ( .A1(c4), .A2(n447), .Z(n443) );
  and2 U352 ( .A1(n450), .A2(n451), .Z(n448) );
  or2 U353 ( .A1(n1999), .A2(n262), .Z(n451) );
  inv1 U354 ( .I(b4), .ZN(n262) );
  or2 U355 ( .A1(b4), .A2(n447), .Z(n450) );
  and2 U356 ( .A1(n452), .A2(n453), .Z(n429) );
  inv1 U357 ( .I(n454), .ZN(n453) );
  and2 U358 ( .A1(n455), .A2(n456), .Z(n454) );
  or2 U359 ( .A1(n456), .A2(n455), .Z(n452) );
  or2 U360 ( .A1(n457), .A2(n458), .Z(n455) );
  and2 U366 ( .A1(n1), .A2(n469), .Z(m7) );
  or2 U367 ( .A1(n470), .A2(n471), .Z(n469) );
  or2 U368 ( .A1(y6), .A2(n472), .Z(n471) );
  and2 U369 ( .A1(e0), .A2(n473), .Z(n472) );
  and2 U370 ( .A1(c0), .A2(g5), .Z(n470) );
  inv1 U371 ( .I(y4), .ZN(m6) );
  inv1 U379 ( .I(n39), .ZN(l9) );
  inv1 U380 ( .I(n29), .ZN(l8) );
  and2 U381 ( .A1(n1), .A2(n480), .Z(l7) );
  or2 U382 ( .A1(n481), .A2(n482), .Z(n480) );
  or2 U383 ( .A1(y6), .A2(n483), .Z(n482) );
  and2 U384 ( .A1(b0), .A2(n473), .Z(n483) );
  and2 U385 ( .A1(g), .A2(g5), .Z(n481) );
  inv1 U386 ( .I(z4), .ZN(l6) );
  inv1 U407 ( .I(n118), .ZN(k9) );
  inv1 U408 ( .I(n46), .ZN(k8) );
  and2 U409 ( .A1(n1), .A2(n507), .Z(k7) );
  or2 U410 ( .A1(n508), .A2(n509), .Z(n507) );
  or2 U411 ( .A1(y6), .A2(n510), .Z(n509) );
  and2 U412 ( .A1(j), .A2(n473), .Z(n510) );
  and2 U413 ( .A1(d0), .A2(g5), .Z(n508) );
  inv1 U414 ( .I(w4), .ZN(k6) );
  or2 U416 ( .A1(n513), .A2(n514), .Z(n512) );
  and2 U417 ( .A1(n1594), .A2(n2022), .Z(n514) );
  or2 U420 ( .A1(n518), .A2(n519), .Z(n517) );
  and2 U422 ( .A1(n519), .A2(n518), .Z(n520) );
  and2 U423 ( .A1(n521), .A2(n522), .Z(n518) );
  inv1 U424 ( .I(n523), .ZN(n522) );
  and2 U425 ( .A1(n524), .A2(n525), .Z(n523) );
  or2 U426 ( .A1(n525), .A2(n524), .Z(n521) );
  or2 U427 ( .A1(n526), .A2(n527), .Z(n524) );
  inv1 U428 ( .I(n528), .ZN(n527) );
  or2 U429 ( .A1(n529), .A2(n530), .Z(n528) );
  and2 U430 ( .A1(n530), .A2(n529), .Z(n526) );
  and2 U431 ( .A1(n531), .A2(n532), .Z(n529) );
  inv1 U432 ( .I(n533), .ZN(n532) );
  and2 U433 ( .A1(n534), .A2(n535), .Z(n533) );
  or2 U434 ( .A1(n535), .A2(n534), .Z(n531) );
  or2 U435 ( .A1(n536), .A2(n537), .Z(n534) );
  and2 U436 ( .A1(n538), .A2(n539), .Z(n537) );
  inv1 U437 ( .I(n540), .ZN(n536) );
  or2 U438 ( .A1(n539), .A2(n538), .Z(n540) );
  inv1 U439 ( .I(n541), .ZN(n538) );
  or2 U440 ( .A1(n542), .A2(n543), .Z(n541) );
  and2 U441 ( .A1(h4), .A2(n544), .Z(n543) );
  or2 U442 ( .A1(n545), .A2(n546), .Z(n544) );
  and2 U443 ( .A1(a3), .A2(v2), .Z(n546) );
  and2 U444 ( .A1(w2), .A2(n216), .Z(n545) );
  and2 U445 ( .A1(n547), .A2(n548), .Z(n542) );
  or2 U446 ( .A1(n549), .A2(n550), .Z(n547) );
  and2 U447 ( .A1(a3), .A2(n551), .Z(n550) );
  and2 U448 ( .A1(n216), .A2(n552), .Z(n549) );
  or2 U449 ( .A1(n553), .A2(n554), .Z(n539) );
  and2 U450 ( .A1(n4), .A2(n555), .Z(n554) );
  or2 U451 ( .A1(n556), .A2(n557), .Z(n555) );
  and2 U452 ( .A1(n2), .A2(v2), .Z(n557) );
  and2 U453 ( .A1(w2), .A2(n239), .Z(n556) );
  and2 U454 ( .A1(n558), .A2(n559), .Z(n553) );
  or2 U455 ( .A1(n560), .A2(n561), .Z(n558) );
  and2 U456 ( .A1(n2), .A2(n551), .Z(n561) );
  and2 U457 ( .A1(n239), .A2(n552), .Z(n560) );
  or2 U458 ( .A1(n562), .A2(n563), .Z(n535) );
  and2 U459 ( .A1(i4), .A2(n564), .Z(n563) );
  or2 U460 ( .A1(n565), .A2(n566), .Z(n564) );
  and2 U461 ( .A1(c3), .A2(v2), .Z(n566) );
  and2 U462 ( .A1(w2), .A2(n221), .Z(n565) );
  and2 U463 ( .A1(n567), .A2(n568), .Z(n562) );
  or2 U464 ( .A1(n569), .A2(n570), .Z(n567) );
  and2 U465 ( .A1(c3), .A2(n551), .Z(n570) );
  and2 U466 ( .A1(n221), .A2(n552), .Z(n569) );
  or2 U467 ( .A1(n571), .A2(n572), .Z(n530) );
  and2 U468 ( .A1(n573), .A2(n574), .Z(n572) );
  inv1 U469 ( .I(n575), .ZN(n571) );
  or2 U470 ( .A1(n574), .A2(n573), .Z(n575) );
  or2 U471 ( .A1(n576), .A2(n577), .Z(n573) );
  and2 U472 ( .A1(n578), .A2(n314), .Z(n577) );
  inv1 U473 ( .I(n579), .ZN(n578) );
  and2 U474 ( .A1(n580), .A2(n579), .Z(n576) );
  or2 U475 ( .A1(n581), .A2(n582), .Z(n579) );
  and2 U476 ( .A1(m4), .A2(n583), .Z(n582) );
  or2 U477 ( .A1(n584), .A2(n585), .Z(n583) );
  and2 U478 ( .A1(l2), .A2(v2), .Z(n585) );
  and2 U479 ( .A1(w2), .A2(n206), .Z(n584) );
  and2 U480 ( .A1(n586), .A2(n2015), .Z(n581) );
  or2 U481 ( .A1(n588), .A2(n589), .Z(n586) );
  and2 U482 ( .A1(l2), .A2(n551), .Z(n589) );
  and2 U483 ( .A1(n206), .A2(n552), .Z(n588) );
  or2 U484 ( .A1(n590), .A2(n591), .Z(n574) );
  and2 U485 ( .A1(p2), .A2(n592), .Z(n591) );
  or2 U486 ( .A1(n593), .A2(n594), .Z(n592) );
  and2 U487 ( .A1(j4), .A2(v2), .Z(n594) );
  and2 U488 ( .A1(n2016), .A2(n551), .Z(n593) );
  and2 U489 ( .A1(n596), .A2(n238), .Z(n590) );
  or2 U490 ( .A1(n597), .A2(n598), .Z(n596) );
  and2 U491 ( .A1(j4), .A2(w2), .Z(n598) );
  and2 U492 ( .A1(n2016), .A2(n552), .Z(n597) );
  or2 U493 ( .A1(n599), .A2(n600), .Z(n525) );
  and2 U494 ( .A1(e4), .A2(n601), .Z(n600) );
  or2 U495 ( .A1(n602), .A2(n603), .Z(n601) );
  and2 U496 ( .A1(e3), .A2(v2), .Z(n603) );
  and2 U497 ( .A1(w2), .A2(n220), .Z(n602) );
  and2 U498 ( .A1(n604), .A2(n605), .Z(n599) );
  or2 U499 ( .A1(n606), .A2(n607), .Z(n604) );
  and2 U500 ( .A1(e3), .A2(n551), .Z(n607) );
  and2 U501 ( .A1(n220), .A2(n552), .Z(n606) );
  or2 U502 ( .A1(n608), .A2(n609), .Z(n519) );
  and2 U503 ( .A1(n610), .A2(n611), .Z(n609) );
  inv1 U504 ( .I(n612), .ZN(n608) );
  or2 U505 ( .A1(n611), .A2(n610), .Z(n612) );
  inv1 U506 ( .I(n613), .ZN(n610) );
  or2 U507 ( .A1(n614), .A2(n615), .Z(n613) );
  and2 U508 ( .A1(r2), .A2(n616), .Z(n615) );
  or2 U509 ( .A1(n617), .A2(n618), .Z(n616) );
  and2 U510 ( .A1(k4), .A2(v2), .Z(n618) );
  and2 U511 ( .A1(n619), .A2(n551), .Z(n617) );
  and2 U512 ( .A1(n620), .A2(n235), .Z(n614) );
  or2 U513 ( .A1(n621), .A2(n622), .Z(n620) );
  and2 U514 ( .A1(k4), .A2(w2), .Z(n622) );
  and2 U515 ( .A1(n619), .A2(n552), .Z(n621) );
  or2 U516 ( .A1(n623), .A2(n624), .Z(n611) );
  and2 U517 ( .A1(y2), .A2(n625), .Z(n624) );
  or2 U518 ( .A1(n626), .A2(n627), .Z(n625) );
  and2 U519 ( .A1(g4), .A2(v2), .Z(n627) );
  and2 U520 ( .A1(n2017), .A2(n551), .Z(n626) );
  and2 U521 ( .A1(n629), .A2(n234), .Z(n623) );
  or2 U522 ( .A1(n630), .A2(n631), .Z(n629) );
  and2 U523 ( .A1(g4), .A2(w2), .Z(n631) );
  and2 U524 ( .A1(n2017), .A2(n552), .Z(n630) );
  and2 U525 ( .A1(u5), .A2(n632), .Z(n513) );
  or2 U526 ( .A1(t5), .A2(w0), .Z(n632) );
  and2 U540 ( .A1(n649), .A2(n1565), .Z(n648) );
  or2 U541 ( .A1(n1565), .A2(n649), .Z(n646) );
  or2 U542 ( .A1(n651), .A2(n652), .Z(n649) );
  and2 U543 ( .A1(n653), .A2(n654), .Z(n652) );
  inv1 U544 ( .I(n655), .ZN(n653) );
  and2 U545 ( .A1(n656), .A2(n655), .Z(n651) );
  or2 U546 ( .A1(n657), .A2(n1992), .Z(n655) );
  and2 U547 ( .A1(n1991), .A2(n660), .Z(n657) );
  inv1 U548 ( .I(n654), .ZN(n656) );
  or2 U549 ( .A1(n189), .A2(n661), .Z(n654) );
  and2 U552 ( .A1(n665), .A2(n660), .Z(n664) );
  or2 U554 ( .A1(n660), .A2(n665), .Z(n666) );
  or2 U555 ( .A1(n667), .A2(n668), .Z(n660) );
  and2 U556 ( .A1(n189), .A2(n669), .Z(n667) );
  and2 U574 ( .A1(n691), .A2(n692), .Z(n189) );
  or2 U604 ( .A1(n727), .A2(n728), .Z(n726) );
  and2 U605 ( .A1(n729), .A2(n2020), .Z(n728) );
  and2 U606 ( .A1(n1983), .A2(n1989), .Z(n727) );
  or2 U626 ( .A1(n755), .A2(n756), .Z(n644) );
  and2 U627 ( .A1(n757), .A2(n758), .Z(n756) );
  inv1 U628 ( .I(n759), .ZN(n755) );
  or2 U629 ( .A1(n758), .A2(n757), .Z(n759) );
  or2 U630 ( .A1(n760), .A2(n761), .Z(n757) );
  and2 U631 ( .A1(n762), .A2(n669), .Z(n761) );
  and2 U632 ( .A1(n763), .A2(n1990), .Z(n760) );
  inv1 U633 ( .I(n765), .ZN(n758) );
  or2 U634 ( .A1(n766), .A2(n767), .Z(n765) );
  and2 U635 ( .A1(n768), .A2(n691), .Z(n767) );
  and2 U636 ( .A1(n769), .A2(n692), .Z(n766) );
  and2 U637 ( .A1(n770), .A2(n771), .Z(n754) );
  inv1 U638 ( .I(n772), .ZN(n771) );
  and2 U639 ( .A1(n773), .A2(n1569), .Z(n772) );
  or2 U640 ( .A1(n1569), .A2(n773), .Z(n770) );
  or2 U641 ( .A1(n775), .A2(n776), .Z(n773) );
  and2 U642 ( .A1(n777), .A2(n668), .Z(n776) );
  inv1 U643 ( .I(n778), .ZN(n777) );
  and2 U644 ( .A1(n779), .A2(n778), .Z(n775) );
  inv1 U645 ( .I(n668), .ZN(n779) );
  or2 U649 ( .A1(n661), .A2(n784), .Z(n783) );
  and2 U650 ( .A1(n784), .A2(n661), .Z(n781) );
  and2 U651 ( .A1(n785), .A2(n786), .Z(j9) );
  or2 U652 ( .A1(n184), .A2(n787), .Z(n786) );
  or2 U653 ( .A1(c8), .A2(n788), .Z(n785) );
  inv1 U654 ( .I(n66), .ZN(j8) );
  and2 U655 ( .A1(n1), .A2(n789), .Z(j7) );
  or2 U656 ( .A1(n790), .A2(n791), .Z(n789) );
  or2 U657 ( .A1(y6), .A2(n792), .Z(n791) );
  and2 U658 ( .A1(h), .A2(n473), .Z(n792) );
  and2 U659 ( .A1(i), .A2(g5), .Z(n790) );
  inv1 U660 ( .I(u2), .ZN(j6) );
  or2 U662 ( .A1(n795), .A2(n796), .Z(n794) );
  and2 U663 ( .A1(n1594), .A2(n504), .Z(n796) );
  and2 U665 ( .A1(n799), .A2(n800), .Z(n798) );
  inv1 U666 ( .I(n801), .ZN(n800) );
  and2 U667 ( .A1(n801), .A2(n802), .Z(n797) );
  inv1 U668 ( .I(n799), .ZN(n802) );
  or2 U669 ( .A1(n803), .A2(n804), .Z(n799) );
  and2 U670 ( .A1(n805), .A2(n806), .Z(n804) );
  inv1 U671 ( .I(n807), .ZN(n806) );
  and2 U672 ( .A1(n807), .A2(n808), .Z(n803) );
  inv1 U673 ( .I(n805), .ZN(n808) );
  or2 U674 ( .A1(n809), .A2(n810), .Z(n805) );
  and2 U675 ( .A1(n811), .A2(n812), .Z(n810) );
  inv1 U676 ( .I(n813), .ZN(n811) );
  and2 U677 ( .A1(n814), .A2(n813), .Z(n809) );
  or2 U678 ( .A1(n815), .A2(n816), .Z(n813) );
  and2 U679 ( .A1(n817), .A2(r4), .Z(n816) );
  and2 U680 ( .A1(n818), .A2(n819), .Z(n817) );
  inv1 U681 ( .I(n820), .ZN(n819) );
  and2 U682 ( .A1(n821), .A2(v2), .Z(n820) );
  or2 U683 ( .A1(v2), .A2(n821), .Z(n818) );
  and2 U684 ( .A1(n822), .A2(n2012), .Z(n815) );
  or2 U685 ( .A1(n824), .A2(n825), .Z(n822) );
  inv1 U686 ( .I(n826), .ZN(n825) );
  or2 U687 ( .A1(n821), .A2(t2), .Z(n826) );
  and2 U688 ( .A1(t2), .A2(n821), .Z(n824) );
  or2 U689 ( .A1(n827), .A2(n828), .Z(n821) );
  and2 U690 ( .A1(q4), .A2(n829), .Z(n828) );
  or2 U691 ( .A1(n830), .A2(n831), .Z(n829) );
  and2 U692 ( .A1(v2), .A2(q3), .Z(n831) );
  and2 U693 ( .A1(w2), .A2(n266), .Z(n830) );
  and2 U694 ( .A1(n832), .A2(n2013), .Z(n827) );
  or2 U695 ( .A1(n834), .A2(n835), .Z(n832) );
  and2 U696 ( .A1(q3), .A2(n551), .Z(n835) );
  and2 U697 ( .A1(n266), .A2(n552), .Z(n834) );
  inv1 U698 ( .I(n812), .ZN(n814) );
  or2 U699 ( .A1(n836), .A2(n837), .Z(n812) );
  and2 U700 ( .A1(x3), .A2(n838), .Z(n837) );
  or2 U701 ( .A1(n839), .A2(n840), .Z(n838) );
  and2 U702 ( .A1(v2), .A2(t4), .Z(n840) );
  and2 U703 ( .A1(n551), .A2(n2011), .Z(n839) );
  and2 U704 ( .A1(n842), .A2(n276), .Z(n836) );
  or2 U705 ( .A1(n843), .A2(n844), .Z(n842) );
  and2 U706 ( .A1(w2), .A2(t4), .Z(n844) );
  and2 U707 ( .A1(n2011), .A2(n552), .Z(n843) );
  or2 U708 ( .A1(n845), .A2(n846), .Z(n807) );
  and2 U709 ( .A1(n847), .A2(n848), .Z(n846) );
  inv1 U710 ( .I(n849), .ZN(n847) );
  and2 U711 ( .A1(n401), .A2(n849), .Z(n845) );
  or2 U712 ( .A1(n850), .A2(n851), .Z(n849) );
  and2 U713 ( .A1(v3), .A2(n852), .Z(n851) );
  or2 U714 ( .A1(n853), .A2(n854), .Z(n852) );
  and2 U715 ( .A1(v2), .A2(s4), .Z(n854) );
  and2 U716 ( .A1(n855), .A2(n551), .Z(n853) );
  and2 U717 ( .A1(n856), .A2(n271), .Z(n850) );
  or2 U718 ( .A1(n857), .A2(n858), .Z(n856) );
  and2 U719 ( .A1(w2), .A2(s4), .Z(n858) );
  and2 U720 ( .A1(n855), .A2(n552), .Z(n857) );
  or2 U721 ( .A1(n859), .A2(n860), .Z(n801) );
  and2 U722 ( .A1(n861), .A2(n862), .Z(n860) );
  inv1 U723 ( .I(n863), .ZN(n862) );
  and2 U724 ( .A1(n863), .A2(n864), .Z(n859) );
  inv1 U725 ( .I(n861), .ZN(n864) );
  or2 U726 ( .A1(n865), .A2(n866), .Z(n861) );
  and2 U727 ( .A1(n867), .A2(n396), .Z(n866) );
  and2 U728 ( .A1(n868), .A2(n400), .Z(n865) );
  or2 U729 ( .A1(n869), .A2(n870), .Z(n863) );
  and2 U730 ( .A1(n871), .A2(n394), .Z(n870) );
  and2 U731 ( .A1(n1986), .A2(n392), .Z(n869) );
  and2 U732 ( .A1(u5), .A2(n873), .Z(n795) );
  or2 U733 ( .A1(t5), .A2(y0), .Z(n873) );
  or2 U741 ( .A1(n882), .A2(n883), .Z(n879) );
  inv1 U742 ( .I(n884), .ZN(n883) );
  or2 U743 ( .A1(n885), .A2(n886), .Z(n884) );
  and2 U744 ( .A1(n886), .A2(n885), .Z(n882) );
  and2 U745 ( .A1(n887), .A2(n888), .Z(n885) );
  inv1 U746 ( .I(n889), .ZN(n888) );
  and2 U747 ( .A1(n1978), .A2(n2018), .Z(n889) );
  or2 U748 ( .A1(n892), .A2(n893), .Z(n886) );
  inv1 U749 ( .I(n894), .ZN(n893) );
  or2 U750 ( .A1(n895), .A2(n896), .Z(n894) );
  and2 U751 ( .A1(n896), .A2(n895), .Z(n892) );
  and2 U752 ( .A1(n2023), .A2(n898), .Z(n895) );
  and2 U757 ( .A1(n2002), .A2(n905), .Z(n902) );
  or2 U760 ( .A1(n909), .A2(n910), .Z(n896) );
  and2 U761 ( .A1(n911), .A2(n447), .Z(n910) );
  inv1 U762 ( .I(n905), .ZN(n911) );
  and2 U763 ( .A1(n1999), .A2(n905), .Z(n909) );
  or2 U764 ( .A1(n912), .A2(n2001), .Z(n905) );
  or2 U780 ( .A1(n933), .A2(n934), .Z(n927) );
  and2 U781 ( .A1(n935), .A2(n2000), .Z(n934) );
  and2 U782 ( .A1(n2024), .A2(n2002), .Z(n933) );
  inv1 U850 ( .I(n1014), .ZN(i9) );
  or2 U851 ( .A1(n1015), .A2(n1016), .Z(n1014) );
  and2 U852 ( .A1(v5), .A2(j1), .Z(n1016) );
  and2 U853 ( .A1(n1017), .A2(n1018), .Z(n1015) );
  or2 U854 ( .A1(o5), .A2(n1019), .Z(n1018) );
  and2 U855 ( .A1(n1020), .A2(n1021), .Z(n1019) );
  or2 U856 ( .A1(n5), .A2(n401), .Z(n1021) );
  inv1 U857 ( .I(n848), .ZN(n401) );
  inv1 U858 ( .I(n1022), .ZN(n1020) );
  and2 U859 ( .A1(b1), .A2(n5), .Z(n1022) );
  or2 U860 ( .A1(n1023), .A2(n1024), .Z(n1017) );
  inv1 U861 ( .I(o5), .ZN(n1024) );
  and2 U862 ( .A1(n1025), .A2(n1026), .Z(n1023) );
  or2 U863 ( .A1(n5), .A2(n788), .Z(n1026) );
  inv1 U864 ( .I(n787), .ZN(n788) );
  or2 U865 ( .A1(n1027), .A2(n1028), .Z(n787) );
  and2 U866 ( .A1(n1985), .A2(n1029), .Z(n1028) );
  inv1 U867 ( .I(i1), .ZN(n1029) );
  and2 U868 ( .A1(i1), .A2(n85), .Z(n1027) );
  inv1 U869 ( .I(n1030), .ZN(n1025) );
  and2 U870 ( .A1(n184), .A2(n5), .Z(n1030) );
  inv1 U871 ( .I(n83), .ZN(i8) );
  or2 U872 ( .A1(y6), .A2(n1031), .Z(i7) );
  inv1 U873 ( .I(f0), .ZN(n1031) );
  inv1 U874 ( .I(n1032), .ZN(y6) );
  and2 U875 ( .A1(o1), .A2(n1), .Z(i6) );
  or2 U876 ( .A1(n1033), .A2(n1034), .Z(i10) );
  or2 U877 ( .A1(n1035), .A2(n1036), .Z(n1034) );
  and2 U878 ( .A1(u1), .A2(n147), .Z(n1036) );
  and2 U879 ( .A1(n148), .A2(n115), .Z(n1035) );
  or2 U880 ( .A1(n1037), .A2(n1038), .Z(n1033) );
  and2 U881 ( .A1(e2), .A2(n152), .Z(n1038) );
  and2 U882 ( .A1(n153), .A2(n118), .Z(n1037) );
  or2 U883 ( .A1(n1039), .A2(n1040), .Z(h9) );
  or2 U884 ( .A1(n1041), .A2(n1042), .Z(n1040) );
  and2 U885 ( .A1(p1), .A2(n147), .Z(n1042) );
  and2 U886 ( .A1(n148), .A2(n66), .Z(n1041) );
  or2 U887 ( .A1(n1043), .A2(n1044), .Z(n1039) );
  and2 U888 ( .A1(q1), .A2(n152), .Z(n1044) );
  and2 U889 ( .A1(n153), .A2(n67), .Z(n1043) );
  or2 U890 ( .A1(n1045), .A2(n1046), .Z(h8) );
  or2 U891 ( .A1(n1047), .A2(n1048), .Z(n1046) );
  and2 U892 ( .A1(v), .A2(n15), .Z(n1048) );
  and2 U893 ( .A1(c), .A2(n16), .Z(n1047) );
  or2 U894 ( .A1(n1049), .A2(n1050), .Z(n1045) );
  and2 U895 ( .A1(n1987), .A2(n149), .Z(n1050) );
  and2 U896 ( .A1(n1997), .A2(n31), .Z(n1049) );
  inv1 U897 ( .I(y3), .ZN(h6) );
  or2 U898 ( .A1(n1051), .A2(n1052), .Z(h10) );
  or2 U899 ( .A1(n1053), .A2(n1054), .Z(n1052) );
  and2 U900 ( .A1(v1), .A2(n147), .Z(n1054) );
  and2 U901 ( .A1(n148), .A2(n38), .Z(n1053) );
  or2 U902 ( .A1(n1055), .A2(n1056), .Z(n1051) );
  and2 U903 ( .A1(f2), .A2(n152), .Z(n1056) );
  and2 U904 ( .A1(n153), .A2(n39), .Z(n1055) );
  or2 U905 ( .A1(n1057), .A2(n1058), .Z(g9) );
  or2 U906 ( .A1(n1059), .A2(n1060), .Z(n1058) );
  and2 U907 ( .A1(r1), .A2(n147), .Z(n1060) );
  and2 U908 ( .A1(n148), .A2(n46), .Z(n1059) );
  or2 U909 ( .A1(n1061), .A2(n1062), .Z(n1057) );
  and2 U910 ( .A1(s1), .A2(n152), .Z(n1062) );
  and2 U911 ( .A1(n153), .A2(n47), .Z(n1061) );
  inv1 U912 ( .I(n47), .ZN(g8) );
  inv1 U913 ( .I(n1063), .ZN(h7) );
  and2 U914 ( .A1(n1064), .A2(n1065), .Z(n1063) );
  or2 U915 ( .A1(m), .A2(n473), .Z(n1065) );
  and2 U916 ( .A1(n1066), .A2(n1032), .Z(n1064) );
  or2 U917 ( .A1(i0), .A2(g5), .Z(n1066) );
  inv1 U918 ( .I(u3), .ZN(g6) );
  or2 U919 ( .A1(n1067), .A2(n1068), .Z(g10) );
  or2 U920 ( .A1(n1069), .A2(n1070), .Z(n1068) );
  and2 U921 ( .A1(w1), .A2(n147), .Z(n1070) );
  and2 U922 ( .A1(n148), .A2(n20), .Z(n1069) );
  or2 U923 ( .A1(n1071), .A2(n1072), .Z(n1067) );
  and2 U924 ( .A1(g2), .A2(n152), .Z(n1072) );
  and2 U925 ( .A1(n153), .A2(n22), .Z(n1071) );
  or2 U926 ( .A1(n1073), .A2(n1074), .Z(f9) );
  or2 U927 ( .A1(n1075), .A2(n1076), .Z(n1074) );
  and2 U928 ( .A1(t1), .A2(n147), .Z(n1076) );
  and2 U929 ( .A1(n148), .A2(n29), .Z(n1075) );
  or2 U930 ( .A1(n1077), .A2(n1078), .Z(n1073) );
  and2 U931 ( .A1(d2), .A2(n152), .Z(n1078) );
  and2 U932 ( .A1(n153), .A2(n30), .Z(n1077) );
  inv1 U933 ( .I(n67), .ZN(f8) );
  inv1 U934 ( .I(n1079), .ZN(f7) );
  and2 U935 ( .A1(n1080), .A2(n1081), .Z(n1079) );
  or2 U936 ( .A1(h0), .A2(n473), .Z(n1081) );
  inv1 U937 ( .I(g5), .ZN(n473) );
  and2 U938 ( .A1(n1082), .A2(n1032), .Z(n1080) );
  and2 U939 ( .A1(k), .A2(l), .Z(n1032) );
  or2 U940 ( .A1(g5), .A2(g0), .Z(n1082) );
  or2 U941 ( .A1(n1083), .A2(n1084), .Z(f10) );
  or2 U942 ( .A1(n1085), .A2(n1086), .Z(n1084) );
  and2 U943 ( .A1(y1), .A2(n147), .Z(n1086) );
  and2 U944 ( .A1(n148), .A2(n54), .Z(n1085) );
  or2 U945 ( .A1(n1087), .A2(n1088), .Z(n1083) );
  and2 U946 ( .A1(i2), .A2(n152), .Z(n1088) );
  and2 U947 ( .A1(n153), .A2(n59), .Z(n1087) );
  or2 U948 ( .A1(n1089), .A2(n1090), .Z(e9) );
  or2 U949 ( .A1(n1091), .A2(n1092), .Z(n1090) );
  and2 U950 ( .A1(x1), .A2(n147), .Z(n1092) );
  and2 U951 ( .A1(n1093), .A2(d5), .Z(n147) );
  and2 U952 ( .A1(n148), .A2(n83), .Z(n1091) );
  and2 U953 ( .A1(n1094), .A2(d5), .Z(n148) );
  or2 U954 ( .A1(n1095), .A2(n1096), .Z(n1089) );
  and2 U955 ( .A1(h2), .A2(n152), .Z(n1096) );
  and2 U956 ( .A1(n2008), .A2(n1093), .Z(n152) );
  and2 U957 ( .A1(l1), .A2(e5), .Z(n1093) );
  and2 U958 ( .A1(n153), .A2(n84), .Z(n1095) );
  and2 U959 ( .A1(n2008), .A2(n1094), .Z(n153) );
  and2 U960 ( .A1(n2007), .A2(l1), .Z(n1094) );
  inv1 U963 ( .I(n84), .ZN(e8) );
  inv1 U964 ( .I(j3), .ZN(e7) );
  or2 U965 ( .A1(n1097), .A2(n1098), .Z(e10) );
  or2 U966 ( .A1(n1099), .A2(n1100), .Z(n1098) );
  and2 U967 ( .A1(u1), .A2(n158), .Z(n1100) );
  and2 U968 ( .A1(n159), .A2(n115), .Z(n1099) );
  or2 U969 ( .A1(n1101), .A2(n1102), .Z(n115) );
  or2 U970 ( .A1(n1103), .A2(n1104), .Z(n1102) );
  and2 U971 ( .A1(n1595), .A2(n296), .Z(n1104) );
  or2 U972 ( .A1(n1105), .A2(n1106), .Z(n296) );
  and2 U973 ( .A1(n1107), .A2(n1108), .Z(n1106) );
  or2 U974 ( .A1(n1109), .A2(n1110), .Z(n1107) );
  and2 U975 ( .A1(n725), .A2(n1111), .Z(n1110) );
  and2 U976 ( .A1(n1112), .A2(n2019), .Z(n1109) );
  inv1 U977 ( .I(n1111), .ZN(n1112) );
  or2 U978 ( .A1(n1979), .A2(n1113), .Z(n1111) );
  and2 U981 ( .A1(n1115), .A2(n1988), .Z(n1105) );
  and2 U982 ( .A1(n1117), .A2(n1118), .Z(n1115) );
  inv1 U983 ( .I(n68), .ZN(n1118) );
  and2 U984 ( .A1(n1113), .A2(n2019), .Z(n68) );
  or2 U985 ( .A1(n2019), .A2(n1113), .Z(n1117) );
  or2 U989 ( .A1(n105), .A2(n1120), .Z(n725) );
  and2 U990 ( .A1(n1980), .A2(n1121), .Z(n1120) );
  and2 U992 ( .A1(l4), .A2(n365), .Z(n105) );
  and2 U994 ( .A1(k2), .A2(t3), .Z(n1123) );
  and2 U996 ( .A1(t0), .A2(n1124), .Z(n1103) );
  and2 U997 ( .A1(n580), .A2(n1594), .Z(n1101) );
  inv1 U998 ( .I(n314), .ZN(n580) );
  or2 U999 ( .A1(n1125), .A2(n1126), .Z(n314) );
  and2 U1000 ( .A1(l4), .A2(n1127), .Z(n1126) );
  or2 U1001 ( .A1(n1128), .A2(n1129), .Z(n1127) );
  and2 U1002 ( .A1(j2), .A2(v2), .Z(n1129) );
  and2 U1003 ( .A1(w2), .A2(n230), .Z(n1128) );
  and2 U1004 ( .A1(n1130), .A2(n1121), .Z(n1125) );
  inv1 U1005 ( .I(l4), .ZN(n1121) );
  or2 U1006 ( .A1(n1131), .A2(n1132), .Z(n1130) );
  and2 U1007 ( .A1(j2), .A2(n551), .Z(n1132) );
  and2 U1008 ( .A1(n230), .A2(n552), .Z(n1131) );
  inv1 U1009 ( .I(j2), .ZN(n230) );
  or2 U1010 ( .A1(n1133), .A2(n1134), .Z(n1097) );
  and2 U1011 ( .A1(e2), .A2(n162), .Z(n1134) );
  and2 U1012 ( .A1(n163), .A2(n118), .Z(n1133) );
  or2 U1013 ( .A1(n1135), .A2(n1136), .Z(n118) );
  or2 U1014 ( .A1(n1137), .A2(n1138), .Z(n1136) );
  and2 U1015 ( .A1(n1595), .A2(n184), .Z(n1138) );
  and2 U1016 ( .A1(b1), .A2(n1124), .Z(n1137) );
  and2 U1017 ( .A1(n1594), .A2(n848), .Z(n1135) );
  or2 U1018 ( .A1(n1139), .A2(n1140), .Z(n848) );
  and2 U1019 ( .A1(t2), .A2(i3), .Z(n1140) );
  and2 U1020 ( .A1(x2), .A2(n267), .Z(n1139) );
  inv1 U1021 ( .I(i3), .ZN(n267) );
  or2 U1022 ( .A1(n1141), .A2(n1142), .Z(d9) );
  or2 U1023 ( .A1(n1143), .A2(n1144), .Z(n1142) );
  and2 U1024 ( .A1(p1), .A2(n158), .Z(n1144) );
  and2 U1025 ( .A1(n159), .A2(n66), .Z(n1143) );
  or2 U1026 ( .A1(n1145), .A2(n1146), .Z(n66) );
  or2 U1027 ( .A1(n1147), .A2(n1148), .Z(n1146) );
  and2 U1028 ( .A1(n1595), .A2(n288), .Z(n1148) );
  or2 U1029 ( .A1(n1149), .A2(n1150), .Z(n288) );
  and2 U1030 ( .A1(n678), .A2(n1151), .Z(n1150) );
  and2 U1031 ( .A1(n1152), .A2(n1991), .Z(n1149) );
  inv1 U1032 ( .I(n1151), .ZN(n1152) );
  and2 U1033 ( .A1(e1), .A2(n1124), .Z(n1147) );
  and2 U1034 ( .A1(n1153), .A2(n1594), .Z(n1145) );
  inv1 U1035 ( .I(n312), .ZN(n1153) );
  or2 U1036 ( .A1(n1154), .A2(n1155), .Z(n312) );
  and2 U1037 ( .A1(y2), .A2(n1156), .Z(n1155) );
  or2 U1038 ( .A1(n1157), .A2(n1158), .Z(n1156) );
  and2 U1039 ( .A1(g4), .A2(n1159), .Z(n1158) );
  and2 U1040 ( .A1(j5), .A2(n2017), .Z(n1157) );
  and2 U1041 ( .A1(n1160), .A2(n234), .Z(n1154) );
  inv1 U1042 ( .I(y2), .ZN(n234) );
  or2 U1043 ( .A1(n1161), .A2(n1162), .Z(n1160) );
  and2 U1044 ( .A1(g4), .A2(n1163), .Z(n1162) );
  and2 U1045 ( .A1(k5), .A2(n2017), .Z(n1161) );
  or2 U1046 ( .A1(n1164), .A2(n1165), .Z(n1141) );
  and2 U1047 ( .A1(q1), .A2(n162), .Z(n1165) );
  and2 U1048 ( .A1(n163), .A2(n67), .Z(n1164) );
  or2 U1049 ( .A1(n1166), .A2(n1167), .Z(n67) );
  or2 U1050 ( .A1(n1168), .A2(n1169), .Z(n1167) );
  and2 U1051 ( .A1(g1), .A2(n1124), .Z(n1169) );
  and2 U1052 ( .A1(n1170), .A2(n1594), .Z(n1168) );
  inv1 U1053 ( .I(n399), .ZN(n1170) );
  or2 U1054 ( .A1(n1171), .A2(n1172), .Z(n399) );
  and2 U1055 ( .A1(r4), .A2(n1159), .Z(n1172) );
  and2 U1056 ( .A1(j5), .A2(n2012), .Z(n1171) );
  and2 U1057 ( .A1(n1595), .A2(n178), .Z(n1166) );
  or2 U1058 ( .A1(n1173), .A2(n1174), .Z(n178) );
  and2 U1059 ( .A1(n935), .A2(n1175), .Z(n1174) );
  and2 U1060 ( .A1(n1176), .A2(n2002), .Z(n1173) );
  inv1 U1061 ( .I(n1175), .ZN(n1176) );
  or2 U1062 ( .A1(n1177), .A2(n1178), .Z(d8) );
  or2 U1063 ( .A1(n1179), .A2(n1180), .Z(n1178) );
  and2 U1064 ( .A1(v), .A2(n52), .Z(n1180) );
  and2 U1065 ( .A1(p5), .A2(q5), .Z(n52) );
  and2 U1066 ( .A1(n53), .A2(n149), .Z(n1179) );
  and2 U1067 ( .A1(n2006), .A2(q5), .Z(n53) );
  or2 U1068 ( .A1(n1182), .A2(n1183), .Z(n1177) );
  and2 U1069 ( .A1(c), .A2(n1981), .Z(n1183) );
  and2 U1071 ( .A1(n1982), .A2(n31), .Z(n1182) );
  or2 U1072 ( .A1(n1185), .A2(n1186), .Z(n31) );
  or2 U1073 ( .A1(n1187), .A2(n1188), .Z(n1186) );
  and2 U1074 ( .A1(n1595), .A2(n180), .Z(n1188) );
  or2 U1075 ( .A1(n1189), .A2(n1190), .Z(n180) );
  and2 U1076 ( .A1(n1999), .A2(n1191), .Z(n1190) );
  and2 U1077 ( .A1(u), .A2(n447), .Z(n1189) );
  and2 U1078 ( .A1(h1), .A2(n1124), .Z(n1187) );
  and2 U1079 ( .A1(n871), .A2(n1594), .Z(n1185) );
  inv1 U1080 ( .I(n392), .ZN(n871) );
  or2 U1081 ( .A1(n1192), .A2(n1193), .Z(n392) );
  and2 U1082 ( .A1(w2), .A2(n275), .Z(n1193) );
  inv1 U1083 ( .I(z3), .ZN(n275) );
  and2 U1084 ( .A1(v2), .A2(z3), .Z(n1192) );
  or2 U1088 ( .A1(n1194), .A2(n1195), .Z(d10) );
  or2 U1089 ( .A1(n1196), .A2(n1197), .Z(n1195) );
  and2 U1090 ( .A1(v1), .A2(n158), .Z(n1197) );
  and2 U1091 ( .A1(n159), .A2(n38), .Z(n1196) );
  or2 U1092 ( .A1(n1198), .A2(n1199), .Z(n38) );
  or2 U1093 ( .A1(n1200), .A2(n1201), .Z(n1199) );
  and2 U1094 ( .A1(n1595), .A2(n298), .Z(n1201) );
  or2 U1095 ( .A1(n1202), .A2(n1203), .Z(n298) );
  and2 U1096 ( .A1(n1204), .A2(n1108), .Z(n1203) );
  or2 U1097 ( .A1(n1205), .A2(n1206), .Z(n1204) );
  and2 U1115 ( .A1(m2), .A2(t3), .Z(n1216) );
  and2 U1120 ( .A1(s0), .A2(n1124), .Z(n1200) );
  and2 U1121 ( .A1(n1219), .A2(n1594), .Z(n1198) );
  inv1 U1122 ( .I(n304), .ZN(n1219) );
  or2 U1123 ( .A1(n1220), .A2(n1221), .Z(n304) );
  and2 U1124 ( .A1(m4), .A2(n1222), .Z(n1221) );
  or2 U1125 ( .A1(n1223), .A2(n1224), .Z(n1222) );
  and2 U1126 ( .A1(l2), .A2(n1159), .Z(n1224) );
  and2 U1127 ( .A1(n206), .A2(n1163), .Z(n1223) );
  and2 U1128 ( .A1(n1225), .A2(n2015), .Z(n1220) );
  or2 U1130 ( .A1(n1226), .A2(n1227), .Z(n1225) );
  and2 U1131 ( .A1(k5), .A2(n206), .Z(n1227) );
  inv1 U1132 ( .I(l2), .ZN(n206) );
  and2 U1133 ( .A1(l2), .A2(j5), .Z(n1226) );
  or2 U1134 ( .A1(n1228), .A2(n1229), .Z(n1194) );
  and2 U1135 ( .A1(f2), .A2(n162), .Z(n1229) );
  and2 U1136 ( .A1(n163), .A2(n39), .Z(n1228) );
  or2 U1137 ( .A1(n1230), .A2(n1231), .Z(n39) );
  or2 U1138 ( .A1(n1232), .A2(n1233), .Z(n1231) );
  and2 U1139 ( .A1(n1595), .A2(n183), .Z(n1233) );
  or2 U1140 ( .A1(n1234), .A2(n1235), .Z(n183) );
  and2 U1151 ( .A1(z0), .A2(n1124), .Z(n1232) );
  and2 U1152 ( .A1(n868), .A2(n1594), .Z(n1230) );
  inv1 U1153 ( .I(n396), .ZN(n868) );
  or2 U1154 ( .A1(n1244), .A2(n1245), .Z(n396) );
  and2 U1155 ( .A1(k3), .A2(v2), .Z(n1245) );
  and2 U1156 ( .A1(w2), .A2(n252), .Z(n1244) );
  inv1 U1157 ( .I(k3), .ZN(n252) );
  or2 U1158 ( .A1(n1246), .A2(n1247), .Z(c9) );
  or2 U1159 ( .A1(n1248), .A2(n1249), .Z(n1247) );
  and2 U1160 ( .A1(r1), .A2(n158), .Z(n1249) );
  and2 U1161 ( .A1(n159), .A2(n46), .Z(n1248) );
  or2 U1162 ( .A1(n1250), .A2(n1251), .Z(n46) );
  or2 U1163 ( .A1(n1252), .A2(n1253), .Z(n1251) );
  and2 U1164 ( .A1(n1595), .A2(n292), .Z(n1253) );
  or2 U1165 ( .A1(n1254), .A2(n1255), .Z(n292) );
  and2 U1166 ( .A1(n763), .A2(n1256), .Z(n1255) );
  inv1 U1167 ( .I(n669), .ZN(n763) );
  and2 U1168 ( .A1(n1257), .A2(n669), .Z(n1254) );
  inv1 U1169 ( .I(n1256), .ZN(n1257) );
  and2 U1170 ( .A1(d1), .A2(n1124), .Z(n1252) );
  and2 U1171 ( .A1(n1258), .A2(n1594), .Z(n1250) );
  inv1 U1172 ( .I(n308), .ZN(n1258) );
  or2 U1173 ( .A1(n1259), .A2(n1260), .Z(n308) );
  and2 U1174 ( .A1(h4), .A2(n1261), .Z(n1260) );
  or2 U1175 ( .A1(n1262), .A2(n1263), .Z(n1261) );
  and2 U1176 ( .A1(a3), .A2(n1159), .Z(n1263) );
  and2 U1177 ( .A1(n216), .A2(n1163), .Z(n1262) );
  and2 U1178 ( .A1(n1264), .A2(n548), .Z(n1259) );
  or2 U1179 ( .A1(n1265), .A2(n1266), .Z(n1264) );
  and2 U1180 ( .A1(j5), .A2(a3), .Z(n1266) );
  and2 U1181 ( .A1(k5), .A2(n216), .Z(n1265) );
  inv1 U1182 ( .I(a3), .ZN(n216) );
  or2 U1183 ( .A1(n1267), .A2(n1268), .Z(n1246) );
  and2 U1184 ( .A1(s1), .A2(n162), .Z(n1268) );
  and2 U1185 ( .A1(n163), .A2(n47), .Z(n1267) );
  or2 U1186 ( .A1(n1269), .A2(n1270), .Z(n47) );
  or2 U1187 ( .A1(n1271), .A2(n1272), .Z(n1270) );
  and2 U1188 ( .A1(n1595), .A2(n179), .Z(n1272) );
  or2 U1189 ( .A1(n1273), .A2(n1274), .Z(n179) );
  and2 U1194 ( .A1(x0), .A2(n1124), .Z(n1271) );
  and2 U1195 ( .A1(n1277), .A2(n1594), .Z(n1269) );
  inv1 U1196 ( .I(n395), .ZN(n1277) );
  or2 U1197 ( .A1(n1278), .A2(n1279), .Z(n395) );
  and2 U1198 ( .A1(v3), .A2(n1280), .Z(n1279) );
  or2 U1199 ( .A1(n1281), .A2(n1282), .Z(n1280) );
  and2 U1200 ( .A1(s4), .A2(n1159), .Z(n1282) );
  and2 U1201 ( .A1(j5), .A2(n855), .Z(n1281) );
  and2 U1202 ( .A1(n1283), .A2(n271), .Z(n1278) );
  inv1 U1203 ( .I(v3), .ZN(n271) );
  or2 U1204 ( .A1(n1284), .A2(n1285), .Z(n1283) );
  and2 U1205 ( .A1(s4), .A2(n1163), .Z(n1285) );
  and2 U1206 ( .A1(k5), .A2(n855), .Z(n1284) );
  inv1 U1207 ( .I(s4), .ZN(n855) );
  inv1 U1208 ( .I(n184), .ZN(c8) );
  or2 U1209 ( .A1(n1286), .A2(n1287), .Z(n184) );
  and2 U1221 ( .A1(s3), .A2(j3), .Z(n1296) );
  and2 U1232 ( .A1(z4), .A2(w4), .Z(c6) );
  or2 U1233 ( .A1(n1302), .A2(n1303), .Z(c10) );
  or2 U1234 ( .A1(n1304), .A2(n1305), .Z(n1303) );
  and2 U1235 ( .A1(w1), .A2(n158), .Z(n1305) );
  and2 U1236 ( .A1(n159), .A2(n20), .Z(n1304) );
  or2 U1237 ( .A1(n1306), .A2(n1307), .Z(n20) );
  or2 U1238 ( .A1(n1308), .A2(n1309), .Z(n1307) );
  and2 U1239 ( .A1(n1595), .A2(n297), .Z(n1309) );
  or2 U1240 ( .A1(n1310), .A2(n1311), .Z(n297) );
  and2 U1241 ( .A1(n1312), .A2(n1108), .Z(n1311) );
  and2 U1247 ( .A1(n1315), .A2(n1988), .Z(n1310) );
  and2 U1261 ( .A1(t), .A2(n1124), .Z(n1308) );
  and2 U1262 ( .A1(n1321), .A2(n1594), .Z(n1306) );
  inv1 U1263 ( .I(n306), .ZN(n1321) );
  or2 U1264 ( .A1(n1322), .A2(n1323), .Z(n306) );
  and2 U1265 ( .A1(n4), .A2(n1324), .Z(n1323) );
  or2 U1266 ( .A1(n1325), .A2(n1326), .Z(n1324) );
  and2 U1267 ( .A1(n2), .A2(n1159), .Z(n1326) );
  and2 U1268 ( .A1(n1163), .A2(n239), .Z(n1325) );
  and2 U1269 ( .A1(n1327), .A2(n559), .Z(n1322) );
  inv1 U1270 ( .I(n4), .ZN(n559) );
  or2 U1271 ( .A1(n1328), .A2(n1329), .Z(n1327) );
  and2 U1272 ( .A1(k5), .A2(n239), .Z(n1329) );
  inv1 U1273 ( .I(n2), .ZN(n239) );
  and2 U1274 ( .A1(j5), .A2(n2), .Z(n1328) );
  or2 U1275 ( .A1(n1330), .A2(n1331), .Z(n1302) );
  and2 U1276 ( .A1(g2), .A2(n162), .Z(n1331) );
  and2 U1277 ( .A1(n163), .A2(n22), .Z(n1330) );
  or2 U1278 ( .A1(n1332), .A2(n1333), .Z(n22) );
  or2 U1279 ( .A1(n1334), .A2(n1335), .Z(n1333) );
  and2 U1280 ( .A1(n1595), .A2(n185), .Z(n1335) );
  or2 U1281 ( .A1(n1336), .A2(n1337), .Z(n185) );
  and2 U1302 ( .A1(u0), .A2(n1124), .Z(n1334) );
  and2 U1303 ( .A1(n1594), .A2(n1986), .Z(n1332) );
  and2 U1306 ( .A1(o4), .A2(n1351), .Z(n1350) );
  or2 U1307 ( .A1(n1352), .A2(n1353), .Z(n1351) );
  and2 U1308 ( .A1(v2), .A2(m3), .Z(n1353) );
  and2 U1309 ( .A1(w2), .A2(n280), .Z(n1352) );
  or2 U1312 ( .A1(n1355), .A2(n1356), .Z(n1354) );
  and2 U1313 ( .A1(m3), .A2(n551), .Z(n1356) );
  and2 U1314 ( .A1(n280), .A2(n552), .Z(n1355) );
  inv1 U1315 ( .I(m3), .ZN(n280) );
  or2 U1316 ( .A1(n1357), .A2(n1358), .Z(b9) );
  or2 U1317 ( .A1(n1359), .A2(n1360), .Z(n1358) );
  and2 U1318 ( .A1(t1), .A2(n158), .Z(n1360) );
  and2 U1319 ( .A1(n159), .A2(n29), .Z(n1359) );
  or2 U1320 ( .A1(n1361), .A2(n1362), .Z(n29) );
  or2 U1321 ( .A1(n1363), .A2(n1364), .Z(n1362) );
  and2 U1322 ( .A1(n1595), .A2(n295), .Z(n1364) );
  or2 U1323 ( .A1(n1365), .A2(n1366), .Z(n295) );
  and2 U1324 ( .A1(n769), .A2(n1367), .Z(n1366) );
  and2 U1325 ( .A1(n1368), .A2(n691), .Z(n1365) );
  inv1 U1326 ( .I(n1367), .ZN(n1368) );
  or2 U1327 ( .A1(n1369), .A2(n784), .Z(n1367) );
  and2 U1328 ( .A1(c1), .A2(n1124), .Z(n1363) );
  and2 U1329 ( .A1(n1370), .A2(n1594), .Z(n1361) );
  inv1 U1330 ( .I(n305), .ZN(n1370) );
  or2 U1331 ( .A1(n1371), .A2(n1372), .Z(n305) );
  and2 U1332 ( .A1(i4), .A2(n1373), .Z(n1372) );
  or2 U1333 ( .A1(n1374), .A2(n1375), .Z(n1373) );
  and2 U1334 ( .A1(c3), .A2(n1159), .Z(n1375) );
  and2 U1335 ( .A1(n221), .A2(n1163), .Z(n1374) );
  and2 U1336 ( .A1(n1376), .A2(n568), .Z(n1371) );
  or2 U1337 ( .A1(n1377), .A2(n1378), .Z(n1376) );
  and2 U1338 ( .A1(j5), .A2(c3), .Z(n1378) );
  and2 U1339 ( .A1(k5), .A2(n221), .Z(n1377) );
  inv1 U1340 ( .I(c3), .ZN(n221) );
  or2 U1341 ( .A1(n1379), .A2(n1380), .Z(n1357) );
  and2 U1342 ( .A1(d2), .A2(n162), .Z(n1380) );
  and2 U1343 ( .A1(n163), .A2(n30), .Z(n1379) );
  inv1 U1344 ( .I(n149), .ZN(b8) );
  or2 U1345 ( .A1(n1381), .A2(n1382), .Z(n149) );
  or2 U1346 ( .A1(n1383), .A2(n1384), .Z(n1382) );
  and2 U1347 ( .A1(n290), .A2(n1595), .Z(n1384) );
  and2 U1348 ( .A1(n1385), .A2(n1386), .Z(n290) );
  or2 U1349 ( .A1(n692), .A2(b), .Z(n1386) );
  or2 U1350 ( .A1(n768), .A2(n1387), .Z(n1385) );
  inv1 U1351 ( .I(b), .ZN(n1387) );
  and2 U1352 ( .A1(v0), .A2(n1124), .Z(n1383) );
  and2 U1353 ( .A1(n1388), .A2(n1594), .Z(n1381) );
  inv1 U1354 ( .I(n313), .ZN(n1388) );
  or2 U1355 ( .A1(n1389), .A2(n1390), .Z(n313) );
  and2 U1356 ( .A1(e4), .A2(n1391), .Z(n1390) );
  or2 U1357 ( .A1(n1392), .A2(n1393), .Z(n1391) );
  and2 U1358 ( .A1(e3), .A2(n1159), .Z(n1393) );
  and2 U1359 ( .A1(n220), .A2(n1163), .Z(n1392) );
  and2 U1360 ( .A1(n1394), .A2(n605), .Z(n1389) );
  or2 U1361 ( .A1(n1395), .A2(n1396), .Z(n1394) );
  and2 U1362 ( .A1(j5), .A2(e3), .Z(n1396) );
  and2 U1363 ( .A1(k5), .A2(n220), .Z(n1395) );
  inv1 U1364 ( .I(e3), .ZN(n220) );
  inv1 U1365 ( .I(a4), .ZN(b6) );
  or2 U1366 ( .A1(n1397), .A2(n1398), .Z(b10) );
  or2 U1367 ( .A1(n1399), .A2(n1400), .Z(n1398) );
  and2 U1368 ( .A1(y1), .A2(n158), .Z(n1400) );
  and2 U1369 ( .A1(n159), .A2(n54), .Z(n1399) );
  or2 U1370 ( .A1(n1401), .A2(n1402), .Z(n1397) );
  and2 U1371 ( .A1(i2), .A2(n162), .Z(n1402) );
  and2 U1372 ( .A1(n163), .A2(n59), .Z(n1401) );
  or2 U1373 ( .A1(n1403), .A2(n1404), .Z(a9) );
  or2 U1374 ( .A1(n1405), .A2(n1406), .Z(n1404) );
  and2 U1375 ( .A1(x1), .A2(n158), .Z(n1406) );
  and2 U1376 ( .A1(n1407), .A2(b5), .Z(n158) );
  and2 U1377 ( .A1(n159), .A2(n83), .Z(n1405) );
  or2 U1378 ( .A1(n1408), .A2(n1409), .Z(n83) );
  or2 U1379 ( .A1(n1410), .A2(n1411), .Z(n1409) );
  and2 U1380 ( .A1(n1595), .A2(n289), .Z(n1411) );
  or2 U1381 ( .A1(n1412), .A2(n1413), .Z(n289) );
  and2 U1382 ( .A1(n762), .A2(n1414), .Z(n1413) );
  and2 U1383 ( .A1(n1415), .A2(n1990), .Z(n1412) );
  inv1 U1384 ( .I(n1414), .ZN(n1415) );
  or2 U1385 ( .A1(n1416), .A2(n1992), .Z(n1414) );
  and2 U1386 ( .A1(n1991), .A2(n1151), .Z(n1416) );
  or2 U1387 ( .A1(n1417), .A2(n1418), .Z(n1151) );
  and2 U1388 ( .A1(n669), .A2(n1256), .Z(n1417) );
  or2 U1389 ( .A1(n1419), .A2(n661), .Z(n1256) );
  and2 U1390 ( .A1(a1), .A2(n1124), .Z(n1410) );
  and2 U1391 ( .A1(n1420), .A2(n1594), .Z(n1408) );
  inv1 U1392 ( .I(n311), .ZN(n1420) );
  or2 U1393 ( .A1(n1421), .A2(n1422), .Z(n311) );
  and2 U1394 ( .A1(r2), .A2(n1423), .Z(n1422) );
  or2 U1395 ( .A1(n1424), .A2(n1425), .Z(n1423) );
  and2 U1396 ( .A1(k4), .A2(n1159), .Z(n1425) );
  and2 U1397 ( .A1(j5), .A2(n619), .Z(n1424) );
  and2 U1398 ( .A1(n1426), .A2(n235), .Z(n1421) );
  inv1 U1399 ( .I(r2), .ZN(n235) );
  or2 U1400 ( .A1(n1427), .A2(n1428), .Z(n1426) );
  and2 U1401 ( .A1(k4), .A2(n1163), .Z(n1428) );
  and2 U1402 ( .A1(k5), .A2(n619), .Z(n1427) );
  and2 U1403 ( .A1(n1429), .A2(b5), .Z(n159) );
  or2 U1404 ( .A1(n1430), .A2(n1431), .Z(n1403) );
  and2 U1405 ( .A1(h2), .A2(n162), .Z(n1431) );
  and2 U1406 ( .A1(n2010), .A2(n1407), .Z(n162) );
  and2 U1407 ( .A1(l1), .A2(c5), .Z(n1407) );
  and2 U1408 ( .A1(n163), .A2(n84), .Z(n1430) );
  or2 U1409 ( .A1(n1432), .A2(n1433), .Z(n84) );
  or2 U1410 ( .A1(n1434), .A2(n1435), .Z(n1433) );
  and2 U1411 ( .A1(n1595), .A2(n177), .Z(n1435) );
  or2 U1412 ( .A1(n1436), .A2(n1437), .Z(n177) );
  and2 U1413 ( .A1(n2003), .A2(n1438), .Z(n1437) );
  and2 U1414 ( .A1(n1439), .A2(n2021), .Z(n1436) );
  inv1 U1415 ( .I(n1438), .ZN(n1439) );
  or2 U1416 ( .A1(n1440), .A2(n903), .Z(n1438) );
  and2 U1417 ( .A1(n2002), .A2(n1175), .Z(n1440) );
  or2 U1418 ( .A1(n1441), .A2(n2001), .Z(n1175) );
  and2 U1422 ( .A1(s), .A2(n1124), .Z(n1434) );
  and2 U1423 ( .A1(n1443), .A2(n1594), .Z(n1432) );
  inv1 U1424 ( .I(n402), .ZN(n1443) );
  or2 U1425 ( .A1(n1444), .A2(n1445), .Z(n402) );
  and2 U1426 ( .A1(q4), .A2(n1446), .Z(n1445) );
  or2 U1427 ( .A1(n1447), .A2(n1448), .Z(n1446) );
  and2 U1428 ( .A1(q3), .A2(n1159), .Z(n1448) );
  and2 U1429 ( .A1(n1163), .A2(n266), .Z(n1447) );
  and2 U1430 ( .A1(n1449), .A2(n2013), .Z(n1444) );
  or2 U1431 ( .A1(n1450), .A2(n1451), .Z(n1449) );
  and2 U1432 ( .A1(k5), .A2(n266), .Z(n1451) );
  inv1 U1433 ( .I(q3), .ZN(n266) );
  and2 U1434 ( .A1(j5), .A2(q3), .Z(n1450) );
  and2 U1435 ( .A1(n2010), .A2(n1429), .Z(n163) );
  and2 U1436 ( .A1(n2009), .A2(l1), .Z(n1429) );
  inv1 U1439 ( .I(n30), .ZN(a8) );
  or2 U1440 ( .A1(n1452), .A2(n1453), .Z(n30) );
  or2 U1441 ( .A1(n1454), .A2(n1455), .Z(n1453) );
  and2 U1442 ( .A1(n1595), .A2(n186), .Z(n1455) );
  inv1 U1445 ( .I(u), .ZN(n1191) );
  and2 U1448 ( .A1(f1), .A2(n1124), .Z(n1454) );
  and2 U1449 ( .A1(n1459), .A2(n1594), .Z(n1452) );
  inv1 U1450 ( .I(n393), .ZN(n1459) );
  or2 U1451 ( .A1(n1460), .A2(n1461), .Z(n393) );
  and2 U1452 ( .A1(x3), .A2(n1462), .Z(n1461) );
  or2 U1453 ( .A1(n1463), .A2(n1464), .Z(n1462) );
  and2 U1454 ( .A1(t4), .A2(n1159), .Z(n1464) );
  and2 U1455 ( .A1(j5), .A2(n2011), .Z(n1463) );
  and2 U1456 ( .A1(n1465), .A2(n276), .Z(n1460) );
  inv1 U1457 ( .I(x3), .ZN(n276) );
  or2 U1458 ( .A1(n1466), .A2(n1467), .Z(n1465) );
  and2 U1459 ( .A1(t4), .A2(n1163), .Z(n1467) );
  and2 U1460 ( .A1(k5), .A2(n2011), .Z(n1466) );
  inv1 U1461 ( .I(w3), .ZN(a6) );
  or2 U1462 ( .A1(n1468), .A2(n1469), .Z(a10) );
  or2 U1463 ( .A1(n1470), .A2(n1471), .Z(n1469) );
  and2 U1464 ( .A1(o), .A2(n15), .Z(n1471) );
  and2 U1465 ( .A1(r5), .A2(s5), .Z(n15) );
  and2 U1466 ( .A1(j0), .A2(n16), .Z(n1470) );
  and2 U1467 ( .A1(n2005), .A2(s5), .Z(n16) );
  or2 U1468 ( .A1(n1473), .A2(n1474), .Z(n1468) );
  and2 U1469 ( .A1(n1987), .A2(n54), .Z(n1474) );
  or2 U1470 ( .A1(n1475), .A2(n1476), .Z(n54) );
  or2 U1471 ( .A1(n1477), .A2(n1478), .Z(n1476) );
  and2 U1472 ( .A1(n1595), .A2(n291), .Z(n1478) );
  or2 U1473 ( .A1(n1479), .A2(n1480), .Z(n291) );
  and2 U1474 ( .A1(n729), .A2(n1108), .Z(n1480) );
  and2 U1475 ( .A1(n1989), .A2(n1988), .Z(n1479) );
  and2 U1481 ( .A1(n1991), .A2(n668), .Z(n1484) );
  or2 U1482 ( .A1(n1485), .A2(n1418), .Z(n668) );
  and2 U1483 ( .A1(n341), .A2(h4), .Z(n1418) );
  and2 U1487 ( .A1(n1419), .A2(n190), .Z(n1481) );
  and2 U1488 ( .A1(n1990), .A2(n1488), .Z(n190) );
  and2 U1489 ( .A1(n669), .A2(n1991), .Z(n1488) );
  and2 U1497 ( .A1(z2), .A2(t3), .Z(n1491) );
  and2 U1499 ( .A1(n1492), .A2(n1493), .Z(n669) );
  or2 U1500 ( .A1(n341), .A2(h4), .Z(n1493) );
  or2 U1501 ( .A1(n548), .A2(n1494), .Z(n1492) );
  and2 U1504 ( .A1(b3), .A2(t3), .Z(n1496) );
  inv1 U1506 ( .I(h4), .ZN(n548) );
  and2 U1509 ( .A1(n1994), .A2(n619), .Z(n1497) );
  inv1 U1510 ( .I(k4), .ZN(n619) );
  and2 U1514 ( .A1(s2), .A2(t3), .Z(n1499) );
  and2 U1516 ( .A1(n1369), .A2(n691), .Z(n1419) );
  inv1 U1517 ( .I(n769), .ZN(n691) );
  or2 U1518 ( .A1(n1487), .A2(n1500), .Z(n769) );
  and2 U1519 ( .A1(n1995), .A2(n568), .Z(n1500) );
  inv1 U1520 ( .I(i4), .ZN(n568) );
  and2 U1522 ( .A1(i4), .A2(n384), .Z(n1487) );
  and2 U1524 ( .A1(d3), .A2(t3), .Z(n1502) );
  and2 U1526 ( .A1(n692), .A2(b), .Z(n1369) );
  inv1 U1527 ( .I(n768), .ZN(n692) );
  or2 U1528 ( .A1(n784), .A2(n665), .Z(n768) );
  and2 U1529 ( .A1(n605), .A2(n1996), .Z(n665) );
  inv1 U1531 ( .I(e4), .ZN(n605) );
  and2 U1532 ( .A1(n380), .A2(e4), .Z(n784) );
  and2 U1534 ( .A1(t3), .A2(f3), .Z(n1504) );
  and2 U1545 ( .A1(r0), .A2(n1124), .Z(n1477) );
  and2 U1546 ( .A1(n1509), .A2(n1594), .Z(n1475) );
  inv1 U1547 ( .I(n307), .ZN(n1509) );
  or2 U1548 ( .A1(n1510), .A2(n1511), .Z(n307) );
  and2 U1549 ( .A1(p2), .A2(n1512), .Z(n1511) );
  or2 U1550 ( .A1(n1513), .A2(n1514), .Z(n1512) );
  and2 U1551 ( .A1(j4), .A2(n1159), .Z(n1514) );
  inv1 U1552 ( .I(m5), .ZN(n1159) );
  and2 U1553 ( .A1(j5), .A2(n2016), .Z(n1513) );
  and2 U1554 ( .A1(n1515), .A2(n238), .Z(n1510) );
  inv1 U1555 ( .I(p2), .ZN(n238) );
  or2 U1556 ( .A1(n1516), .A2(n1517), .Z(n1515) );
  and2 U1557 ( .A1(j4), .A2(n1163), .Z(n1517) );
  inv1 U1558 ( .I(l5), .ZN(n1163) );
  and2 U1559 ( .A1(k5), .A2(n2016), .Z(n1516) );
  and2 U1562 ( .A1(n1997), .A2(n59), .Z(n1473) );
  or2 U1563 ( .A1(n1519), .A2(n1520), .Z(n59) );
  or2 U1564 ( .A1(n1521), .A2(n1522), .Z(n1520) );
  and2 U1565 ( .A1(n1595), .A2(n1998), .Z(n1522) );
  and2 U1591 ( .A1(r3), .A2(s3), .Z(n1536) );
  and2 U1620 ( .A1(s3), .A2(w3), .Z(n1546) );
  and2 U1631 ( .A1(q0), .A2(n1124), .Z(n1521) );
  and2 U1632 ( .A1(n2004), .A2(u5), .Z(n1124) );
  and2 U1633 ( .A1(n867), .A2(n1594), .Z(n1519) );
  inv1 U1637 ( .I(n400), .ZN(n867) );
  or2 U1638 ( .A1(n1553), .A2(n1554), .Z(n400) );
  and2 U1639 ( .A1(p4), .A2(n1555), .Z(n1554) );
  or2 U1640 ( .A1(n1556), .A2(n1557), .Z(n1555) );
  and2 U1641 ( .A1(v2), .A2(o3), .Z(n1557) );
  and2 U1642 ( .A1(w2), .A2(n279), .Z(n1556) );
  and2 U1643 ( .A1(n1558), .A2(n2014), .Z(n1553) );
  or2 U1645 ( .A1(n1559), .A2(n1560), .Z(n1558) );
  and2 U1646 ( .A1(o3), .A2(n551), .Z(n1560) );
  inv1 U1647 ( .I(t2), .ZN(n551) );
  and2 U1648 ( .A1(n279), .A2(n552), .Z(n1559) );
  inv1 U1649 ( .I(x2), .ZN(n552) );
  inv1 U1650 ( .I(o3), .ZN(n279) );
  and2 U1657 ( .A1(n1858), .A2(n1859), .Z(n1564) );
  inv1 U1658 ( .I(n1564), .ZN(n1861) );
  and2 U1659 ( .A1(n666), .A2(n1566), .Z(n1565) );
  inv1 U1660 ( .I(n664), .ZN(n1566) );
  and2 U1661 ( .A1(n1862), .A2(n1860), .Z(n1567) );
  inv1 U1662 ( .I(n1567), .ZN(n1856) );
  and2 U1664 ( .A1(n1570), .A2(n783), .Z(n1569) );
  inv1 U1665 ( .I(n781), .ZN(n1570) );
  inv1 U1667 ( .I(n1571), .ZN(n1875) );
  inv1 U1668 ( .I(n1690), .ZN(n1572) );
  inv1 U1671 ( .I(n1574), .ZN(n1880) );
  or2 U1674 ( .A1(n1948), .A2(n1595), .Z(n1576) );
  or2 U1675 ( .A1(n1946), .A2(n1948), .Z(n1577) );
  and2 U1676 ( .A1(n1801), .A2(n1580), .Z(n1578) );
  or2 U1677 ( .A1(n1578), .A2(n1579), .Z(n1806) );
  and2 U1678 ( .A1(n1985), .A2(n1803), .Z(n1579) );
  and2 U1679 ( .A1(n1984), .A2(n1985), .Z(n1580) );
  inv1 U1682 ( .I(n1568), .ZN(n1766) );
  or2 U1683 ( .A1(n1973), .A2(n1586), .Z(n1584) );
  and2 U1684 ( .A1(n1584), .A2(n1585), .Z(o10) );
  or2 U1685 ( .A1(n1976), .A2(n1975), .Z(n1585) );
  or2 U1686 ( .A1(e5), .A2(n1976), .Z(n1586) );
  or2 U1687 ( .A1(n1810), .A2(n1806), .Z(n1587) );
  or2 U1690 ( .A1(n1666), .A2(n1665), .Z(n1590) );
  inv1 U1694 ( .I(n1592), .ZN(n1801) );
  inv1 U1695 ( .I(n1800), .ZN(n1593) );
  inv1 U1696 ( .I(n1939), .ZN(n1594) );
  inv1 U1697 ( .I(n1932), .ZN(n1595) );
  inv1 U1698 ( .I(p4), .ZN(n2014) );
  or2 U1699 ( .A1(t5), .A2(u5), .Z(n1939) );
  inv1 U1700 ( .I(t5), .ZN(n2004) );
  or2 U1701 ( .A1(n2004), .A2(u5), .Z(n1932) );
  and2 U1703 ( .A1(q3), .A2(n1722), .Z(n1596) );
  or2 U1704 ( .A1(n1596), .A2(n1536), .Z(n1721) );
  inv1 U1705 ( .I(n1721), .ZN(n1719) );
  and2 U1706 ( .A1(q4), .A2(n1719), .Z(n1598) );
  inv1 U1707 ( .I(q4), .ZN(n2013) );
  and2 U1708 ( .A1(n2013), .A2(n1721), .Z(n1597) );
  or2 U1709 ( .A1(n1598), .A2(n1597), .Z(n2021) );
  inv1 U1710 ( .I(r4), .ZN(n2012) );
  or2 U1711 ( .A1(n1722), .A2(u3), .Z(n1718) );
  inv1 U1712 ( .I(n1718), .ZN(n1720) );
  and2 U1713 ( .A1(n2012), .A2(n1720), .Z(n1599) );
  or2 U1714 ( .A1(n1720), .A2(n2012), .Z(n1706) );
  inv1 U1715 ( .I(n1706), .ZN(n903) );
  or2 U1716 ( .A1(n1599), .A2(n903), .Z(n935) );
  and2 U1717 ( .A1(v3), .A2(n1722), .Z(n1600) );
  or2 U1718 ( .A1(n1600), .A2(n1546), .Z(n456) );
  inv1 U1719 ( .I(n456), .ZN(n1601) );
  and2 U1720 ( .A1(n855), .A2(n1601), .Z(n1603) );
  or2 U1721 ( .A1(n1601), .A2(n855), .Z(n1602) );
  inv1 U1722 ( .I(n1602), .ZN(n2001) );
  or2 U1723 ( .A1(n1603), .A2(n2001), .Z(n2024) );
  and2 U1724 ( .A1(a4), .A2(s3), .Z(n1605) );
  and2 U1725 ( .A1(z3), .A2(n1722), .Z(n1604) );
  or2 U1726 ( .A1(n1605), .A2(n1604), .Z(n447) );
  and2 U1727 ( .A1(p3), .A2(s3), .Z(n1607) );
  or2 U1730 ( .A1(n1731), .A2(p4), .Z(n1649) );
  inv1 U1731 ( .I(n1649), .ZN(n1808) );
  inv1 U1734 ( .I(n1780), .ZN(n1779) );
  inv1 U1736 ( .I(t4), .ZN(n2011) );
  and2 U1737 ( .A1(y3), .A2(s3), .Z(n1609) );
  or2 U1739 ( .A1(n1609), .A2(n1608), .Z(n1725) );
  inv1 U1740 ( .I(n1725), .ZN(n1724) );
  and2 U1741 ( .A1(n2011), .A2(n1724), .Z(n1611) );
  or2 U1742 ( .A1(n1724), .A2(n2011), .Z(n1610) );
  inv1 U1743 ( .I(n1610), .ZN(n1703) );
  or2 U1744 ( .A1(n1611), .A2(n1703), .Z(n1712) );
  or2 U1745 ( .A1(n1712), .A2(n447), .Z(n1637) );
  inv1 U1746 ( .I(n2021), .ZN(n2003) );
  or2 U1747 ( .A1(n1637), .A2(n2003), .Z(n1613) );
  or2 U1748 ( .A1(n935), .A2(n2024), .Z(n1612) );
  or2 U1749 ( .A1(n1613), .A2(n1612), .Z(n1747) );
  inv1 U1750 ( .I(n1747), .ZN(n1784) );
  and2 U1751 ( .A1(u), .A2(n1784), .Z(n1619) );
  and2 U1752 ( .A1(q4), .A2(n1721), .Z(n1618) );
  inv1 U1753 ( .I(n935), .ZN(n2002) );
  inv1 U1754 ( .I(n2024), .ZN(n2000) );
  inv1 U1755 ( .I(n1712), .ZN(n1713) );
  and2 U1758 ( .A1(n2000), .A2(n1820), .Z(n1615) );
  or2 U1759 ( .A1(n1615), .A2(n2001), .Z(n1825) );
  and2 U1760 ( .A1(n2002), .A2(n1825), .Z(n1616) );
  or2 U1761 ( .A1(n1616), .A2(n903), .Z(n1759) );
  and2 U1762 ( .A1(n2021), .A2(n1759), .Z(n1617) );
  or2 U1763 ( .A1(n1618), .A2(n1617), .Z(n1785) );
  or2 U1764 ( .A1(n1619), .A2(n1785), .Z(n1685) );
  inv1 U1765 ( .I(n1685), .ZN(n1677) );
  and2 U1766 ( .A1(n1663), .A2(n1677), .Z(n1621) );
  inv1 U1767 ( .I(n1663), .ZN(n1809) );
  and2 U1768 ( .A1(n1809), .A2(n1685), .Z(n1620) );
  or2 U1769 ( .A1(n1621), .A2(n1620), .Z(n1622) );
  inv1 U1770 ( .I(n1622), .ZN(n1998) );
  or2 U1771 ( .A1(r5), .A2(s5), .Z(n1623) );
  inv1 U1772 ( .I(n1623), .ZN(n1997) );
  inv1 U1773 ( .I(j4), .ZN(n2016) );
  and2 U1775 ( .A1(e3), .A2(n1734), .Z(n1624) );
  or2 U1776 ( .A1(n1624), .A2(n1504), .Z(n380) );
  inv1 U1777 ( .I(n380), .ZN(n1996) );
  or2 U1779 ( .A1(n1625), .A2(n1502), .Z(n384) );
  inv1 U1780 ( .I(n384), .ZN(n1995) );
  and2 U1781 ( .A1(r2), .A2(n1734), .Z(n1626) );
  or2 U1782 ( .A1(n1626), .A2(n1499), .Z(n378) );
  inv1 U1783 ( .I(n378), .ZN(n1994) );
  and2 U1784 ( .A1(a3), .A2(n1734), .Z(n1627) );
  or2 U1785 ( .A1(n1627), .A2(n1496), .Z(n341) );
  inv1 U1786 ( .I(n341), .ZN(n1494) );
  and2 U1787 ( .A1(y2), .A2(n1734), .Z(n1628) );
  or2 U1788 ( .A1(n1628), .A2(n1491), .Z(n386) );
  inv1 U1789 ( .I(n386), .ZN(n1993) );
  inv1 U1790 ( .I(g4), .ZN(n2017) );
  or2 U1791 ( .A1(n1993), .A2(n2017), .Z(n1629) );
  inv1 U1792 ( .I(n1629), .ZN(n1992) );
  and2 U1793 ( .A1(n2017), .A2(n1993), .Z(n1630) );
  or2 U1794 ( .A1(n1992), .A2(n1630), .Z(n678) );
  inv1 U1795 ( .I(n678), .ZN(n1991) );
  or2 U1796 ( .A1(n1994), .A2(n619), .Z(n1631) );
  inv1 U1797 ( .I(n1631), .ZN(n1634) );
  or2 U1798 ( .A1(n1634), .A2(n1497), .Z(n762) );
  inv1 U1799 ( .I(n762), .ZN(n1990) );
  and2 U1800 ( .A1(q2), .A2(t3), .Z(n1633) );
  or2 U1802 ( .A1(n1633), .A2(n1632), .Z(n1739) );
  or2 U1803 ( .A1(n1739), .A2(j4), .Z(n1854) );
  inv1 U1804 ( .I(n1854), .ZN(n1852) );
  inv1 U1805 ( .I(n1739), .ZN(n1737) );
  or2 U1806 ( .A1(n1737), .A2(n2016), .Z(n1887) );
  or2 U1810 ( .A1(n1992), .A2(n1484), .Z(n778) );
  and2 U1811 ( .A1(n778), .A2(n1990), .Z(n1635) );
  or2 U1812 ( .A1(n1635), .A2(n1634), .Z(n109) );
  or2 U1813 ( .A1(n109), .A2(n1481), .Z(n1108) );
  inv1 U1814 ( .I(n1108), .ZN(n1988) );
  inv1 U1815 ( .I(r5), .ZN(n2005) );
  or2 U1816 ( .A1(n2005), .A2(s5), .Z(n1957) );
  inv1 U1817 ( .I(n1957), .ZN(n1987) );
  or2 U1818 ( .A1(n447), .A2(u), .Z(n1636) );
  and2 U1819 ( .A1(n1712), .A2(n1636), .Z(n1639) );
  inv1 U1820 ( .I(n1637), .ZN(n1705) );
  and2 U1821 ( .A1(n1191), .A2(n1705), .Z(n1638) );
  or2 U1822 ( .A1(n1639), .A2(n1638), .Z(n186) );
  inv1 U1823 ( .I(c5), .ZN(n2009) );
  inv1 U1824 ( .I(b5), .ZN(n2010) );
  and2 U1825 ( .A1(u), .A2(n1713), .Z(n1640) );
  or2 U1826 ( .A1(n1640), .A2(n1820), .Z(n1675) );
  and2 U1827 ( .A1(n2000), .A2(n1675), .Z(n1441) );
  inv1 U1828 ( .I(o4), .ZN(n1644) );
  and2 U1829 ( .A1(n1354), .A2(n1644), .Z(n1641) );
  or2 U1830 ( .A1(n1641), .A2(n1350), .Z(n394) );
  inv1 U1831 ( .I(n394), .ZN(n1986) );
  and2 U1833 ( .A1(n3), .A2(s3), .Z(n1642) );
  inv1 U1835 ( .I(n1728), .ZN(n1730) );
  and2 U1837 ( .A1(n1644), .A2(n1728), .Z(n1645) );
  or2 U1840 ( .A1(n1799), .A2(n1780), .Z(n1664) );
  and2 U1841 ( .A1(n1677), .A2(n1664), .Z(n1648) );
  or2 U1842 ( .A1(n1764), .A2(n1779), .Z(n1647) );
  and2 U1843 ( .A1(n1648), .A2(n1647), .Z(n1336) );
  and2 U1844 ( .A1(n1649), .A2(n1799), .Z(n1651) );
  and2 U1845 ( .A1(n1808), .A2(n1764), .Z(n1650) );
  or2 U1846 ( .A1(n1651), .A2(n1650), .Z(n1652) );
  and2 U1847 ( .A1(n1685), .A2(n1652), .Z(n1337) );
  and2 U1848 ( .A1(o2), .A2(t3), .Z(n1654) );
  or2 U1850 ( .A1(n1654), .A2(n1653), .Z(n1742) );
  inv1 U1851 ( .I(n1742), .ZN(n1744) );
  and2 U1852 ( .A1(n4), .A2(n1744), .Z(n1656) );
  and2 U1853 ( .A1(n559), .A2(n1742), .Z(n1655) );
  or2 U1855 ( .A1(n1880), .A2(n1884), .Z(n1657) );
  and2 U1856 ( .A1(n1689), .A2(n1657), .Z(n1315) );
  and2 U1857 ( .A1(n1852), .A2(n1880), .Z(n1659) );
  and2 U1858 ( .A1(n1854), .A2(n1574), .Z(n1658) );
  or2 U1859 ( .A1(n1659), .A2(n1658), .Z(n1312) );
  and2 U1860 ( .A1(i3), .A2(n1722), .Z(n1660) );
  or2 U1861 ( .A1(n1660), .A2(n1296), .Z(n85) );
  and2 U1862 ( .A1(l3), .A2(s3), .Z(n1662) );
  and2 U1863 ( .A1(k3), .A2(n1722), .Z(n1661) );
  or2 U1864 ( .A1(n1662), .A2(n1661), .Z(n425) );
  and2 U1866 ( .A1(o4), .A2(n1728), .Z(n1665) );
  or2 U1870 ( .A1(n1795), .A2(n85), .Z(n1667) );
  and2 U1871 ( .A1(n1685), .A2(n1667), .Z(n1670) );
  inv1 U1872 ( .I(n85), .ZN(n1985) );
  or2 U1873 ( .A1(n1668), .A2(n1985), .Z(n1669) );
  and2 U1874 ( .A1(n1670), .A2(n1669), .Z(n1286) );
  inv1 U1875 ( .I(n1753), .ZN(n1765) );
  or2 U1876 ( .A1(n1765), .A2(n85), .Z(n1671) );
  and2 U1877 ( .A1(n1677), .A2(n1671), .Z(n1673) );
  or2 U1878 ( .A1(n1753), .A2(n1985), .Z(n1672) );
  and2 U1879 ( .A1(n1673), .A2(n1672), .Z(n1287) );
  inv1 U1880 ( .I(n1675), .ZN(n1674) );
  and2 U1881 ( .A1(n2000), .A2(n1674), .Z(n1273) );
  and2 U1882 ( .A1(n2024), .A2(n1675), .Z(n1274) );
  inv1 U1883 ( .I(n1794), .ZN(n1680) );
  or2 U1884 ( .A1(n1680), .A2(n425), .Z(n1676) );
  and2 U1885 ( .A1(n1677), .A2(n1676), .Z(n1679) );
  inv1 U1886 ( .I(n425), .ZN(n1984) );
  or2 U1887 ( .A1(n1794), .A2(n1984), .Z(n1678) );
  and2 U1888 ( .A1(n1679), .A2(n1678), .Z(n1234) );
  and2 U1889 ( .A1(n1680), .A2(n1766), .Z(n1681) );
  or2 U1890 ( .A1(n1681), .A2(n1984), .Z(n1682) );
  inv1 U1891 ( .I(n1682), .ZN(n1683) );
  or2 U1892 ( .A1(n1683), .A2(n1795), .Z(n1684) );
  and2 U1893 ( .A1(n1685), .A2(n1684), .Z(n1235) );
  inv1 U1894 ( .I(m4), .ZN(n2015) );
  or2 U1896 ( .A1(n1686), .A2(n1216), .Z(n1736) );
  inv1 U1897 ( .I(n1736), .ZN(n1738) );
  and2 U1898 ( .A1(m4), .A2(n1738), .Z(n1688) );
  and2 U1899 ( .A1(n2015), .A2(n1736), .Z(n1687) );
  or2 U1900 ( .A1(n1688), .A2(n1687), .Z(n2020) );
  and2 U1901 ( .A1(n1989), .A2(n1880), .Z(n1691) );
  and2 U1902 ( .A1(n4), .A2(n1742), .Z(n1690) );
  or2 U1903 ( .A1(n1691), .A2(n1875), .Z(n1853) );
  inv1 U1904 ( .I(n1853), .ZN(n1855) );
  and2 U1905 ( .A1(n2020), .A2(n1855), .Z(n1205) );
  or2 U1906 ( .A1(n1855), .A2(n2020), .Z(n1692) );
  inv1 U1907 ( .I(n1692), .ZN(n1206) );
  inv1 U1908 ( .I(n2020), .ZN(n1983) );
  or2 U1909 ( .A1(n1875), .A2(n1983), .Z(n1694) );
  or2 U1910 ( .A1(n1571), .A2(n2020), .Z(n1693) );
  and2 U1911 ( .A1(n1694), .A2(n1693), .Z(n1695) );
  or2 U1912 ( .A1(n1695), .A2(n1108), .Z(n1696) );
  inv1 U1913 ( .I(n1696), .ZN(n1202) );
  inv1 U1914 ( .I(n447), .ZN(n1999) );
  or2 U1915 ( .A1(p5), .A2(q5), .Z(n1697) );
  inv1 U1916 ( .I(n1697), .ZN(n1982) );
  inv1 U1917 ( .I(p5), .ZN(n2006) );
  or2 U1918 ( .A1(n2006), .A2(q5), .Z(n1698) );
  inv1 U1919 ( .I(n1698), .ZN(n1981) );
  and2 U1920 ( .A1(j2), .A2(n1734), .Z(n1699) );
  or2 U1921 ( .A1(n1699), .A2(n1123), .Z(n365) );
  inv1 U1922 ( .I(n365), .ZN(n1980) );
  inv1 U1923 ( .I(n725), .ZN(n2019) );
  or2 U1925 ( .A1(n1738), .A2(n2015), .Z(n1700) );
  inv1 U1927 ( .I(n1876), .ZN(n1113) );
  or2 U1928 ( .A1(n729), .A2(n1983), .Z(n1702) );
  or2 U1929 ( .A1(n1702), .A2(n1574), .Z(n1849) );
  inv1 U1930 ( .I(n1849), .ZN(n1979) );
  inv1 U1931 ( .I(e5), .ZN(n2007) );
  inv1 U1932 ( .I(d5), .ZN(n2008) );
  or2 U1933 ( .A1(n1713), .A2(n1703), .Z(n1704) );
  and2 U1934 ( .A1(n2000), .A2(n1704), .Z(n912) );
  or2 U1935 ( .A1(n1705), .A2(n1820), .Z(n1709) );
  inv1 U1936 ( .I(n902), .ZN(n1707) );
  and2 U1937 ( .A1(n1707), .A2(n1706), .Z(n1708) );
  or2 U1938 ( .A1(n1709), .A2(n1708), .Z(n2023) );
  inv1 U1939 ( .I(n1709), .ZN(n1710) );
  or2 U1940 ( .A1(n1710), .A2(n903), .Z(n1711) );
  or2 U1941 ( .A1(n1711), .A2(n902), .Z(n898) );
  and2 U1942 ( .A1(n2003), .A2(n1712), .Z(n1715) );
  and2 U1943 ( .A1(n2021), .A2(n1713), .Z(n1714) );
  or2 U1944 ( .A1(n1715), .A2(n1714), .Z(n1716) );
  inv1 U1945 ( .I(n1716), .ZN(n1978) );
  inv1 U1946 ( .I(n927), .ZN(n2018) );
  or2 U1947 ( .A1(n1978), .A2(n2018), .Z(n887) );
  or2 U1948 ( .A1(n798), .A2(n797), .Z(n504) );
  inv1 U1949 ( .I(n517), .ZN(n1717) );
  or2 U1950 ( .A1(n520), .A2(n1717), .Z(n2022) );
  and2 U1951 ( .A1(n1719), .A2(n1718), .Z(n457) );
  and2 U1952 ( .A1(n1721), .A2(n1720), .Z(n458) );
  and2 U1953 ( .A1(n448), .A2(n1722), .Z(n1723) );
  or2 U1954 ( .A1(n1723), .A2(n441), .Z(n434) );
  and2 U1955 ( .A1(n85), .A2(n1724), .Z(n1727) );
  and2 U1956 ( .A1(n1985), .A2(n1725), .Z(n1726) );
  or2 U1957 ( .A1(n1727), .A2(n1726), .Z(n433) );
  and2 U1958 ( .A1(n1729), .A2(n1728), .Z(n1733) );
  and2 U1959 ( .A1(n1731), .A2(n1730), .Z(n1732) );
  or2 U1960 ( .A1(n1733), .A2(n1732), .Z(n420) );
  and2 U1961 ( .A1(n366), .A2(n1734), .Z(n1735) );
  or2 U1962 ( .A1(n1735), .A2(n359), .Z(n350) );
  and2 U1963 ( .A1(n1737), .A2(n1736), .Z(n1741) );
  and2 U1964 ( .A1(n1739), .A2(n1738), .Z(n1740) );
  or2 U1965 ( .A1(n1741), .A2(n1740), .Z(n349) );
  inv1 U1966 ( .I(n373), .ZN(n1743) );
  and2 U1967 ( .A1(n1743), .A2(n1742), .Z(n1746) );
  and2 U1968 ( .A1(n373), .A2(n1744), .Z(n1745) );
  or2 U1969 ( .A1(n1746), .A2(n1745), .Z(n345) );
  or2 U1970 ( .A1(n1747), .A2(n85), .Z(n1749) );
  or2 U1971 ( .A1(n1766), .A2(n425), .Z(n1748) );
  or2 U1972 ( .A1(n1749), .A2(n1748), .Z(n1750) );
  inv1 U1973 ( .I(n1750), .ZN(q7) );
  or2 U1974 ( .A1(n1876), .A2(n725), .Z(n1751) );
  inv1 U1975 ( .I(n1751), .ZN(n1752) );
  or2 U1976 ( .A1(n1752), .A2(n69), .Z(v7) );
  or2 U1977 ( .A1(n1753), .A2(n85), .Z(n1755) );
  and2 U1978 ( .A1(n1785), .A2(n1568), .Z(n1754) );
  or2 U1979 ( .A1(n1755), .A2(n1754), .Z(y7) );
  and2 U1980 ( .A1(n2018), .A2(n1978), .Z(n1757) );
  inv1 U1981 ( .I(n887), .ZN(n1756) );
  or2 U1982 ( .A1(n1757), .A2(n1756), .Z(n1760) );
  inv1 U1983 ( .I(n1760), .ZN(n1758) );
  and2 U1984 ( .A1(n1759), .A2(n1758), .Z(n1763) );
  inv1 U1985 ( .I(n1759), .ZN(n1761) );
  and2 U1986 ( .A1(n1761), .A2(n1760), .Z(n1762) );
  or2 U1987 ( .A1(n1763), .A2(n1762), .Z(n1831) );
  or2 U1988 ( .A1(n1764), .A2(n1809), .Z(n1769) );
  or2 U1989 ( .A1(n1765), .A2(n1794), .Z(n1768) );
  and2 U1990 ( .A1(n1766), .A2(n1768), .Z(n1767) );
  and2 U1991 ( .A1(n1769), .A2(n1767), .Z(n1774) );
  inv1 U1992 ( .I(n1768), .ZN(n1772) );
  inv1 U1993 ( .I(n1769), .ZN(n1770) );
  or2 U1994 ( .A1(n1770), .A2(n1568), .Z(n1771) );
  and2 U1995 ( .A1(n1772), .A2(n1771), .Z(n1773) );
  or2 U1996 ( .A1(n1774), .A2(n1773), .Z(n1776) );
  inv1 U1997 ( .I(n1776), .ZN(n1775) );
  and2 U1998 ( .A1(n425), .A2(n1775), .Z(n1778) );
  and2 U1999 ( .A1(n1984), .A2(n1776), .Z(n1777) );
  or2 U2000 ( .A1(n1778), .A2(n1777), .Z(n1789) );
  and2 U2001 ( .A1(n85), .A2(n1779), .Z(n1782) );
  and2 U2002 ( .A1(n1985), .A2(n1780), .Z(n1781) );
  or2 U2003 ( .A1(n1782), .A2(n1781), .Z(n1790) );
  inv1 U2004 ( .I(n1790), .ZN(n1783) );
  or2 U2005 ( .A1(n1789), .A2(n1783), .Z(n1788) );
  and2 U2006 ( .A1(f5), .A2(n1784), .Z(n1786) );
  or2 U2007 ( .A1(n1786), .A2(n1785), .Z(n1812) );
  inv1 U2008 ( .I(n1812), .ZN(n1787) );
  inv1 U2010 ( .I(n1789), .ZN(n1791) );
  or2 U2011 ( .A1(n1791), .A2(n1790), .Z(n1792) );
  or2 U2013 ( .A1(n1795), .A2(n1590), .Z(n1798) );
  or2 U2014 ( .A1(n1798), .A2(n1799), .Z(n1796) );
  and2 U2016 ( .A1(n1799), .A2(n1798), .Z(n1800) );
  and2 U2018 ( .A1(n1984), .A2(n1801), .Z(n1802) );
  or2 U2019 ( .A1(n1803), .A2(n1802), .Z(n1805) );
  or2 U2022 ( .A1(n1807), .A2(n1806), .Z(n1813) );
  or2 U2023 ( .A1(n1809), .A2(n1808), .Z(n1814) );
  inv1 U2024 ( .I(n1814), .ZN(n1810) );
  or2 U2025 ( .A1(n1587), .A2(n1807), .Z(n1811) );
  inv1 U2027 ( .I(n1813), .ZN(n1815) );
  inv1 U2033 ( .I(n1820), .ZN(n1821) );
  and2 U2034 ( .A1(n1589), .A2(n1821), .Z(n1822) );
  inv1 U2036 ( .I(n1827), .ZN(n1824) );
  inv1 U2038 ( .I(n1825), .ZN(n1826) );
  and2 U2039 ( .A1(n1827), .A2(n1826), .Z(n1828) );
  inv1 U2041 ( .I(n1833), .ZN(n1830) );
  inv1 U2043 ( .I(n1831), .ZN(n1832) );
  or2 U2046 ( .A1(n1943), .A2(f5), .Z(n1836) );
  inv1 U2047 ( .I(n1836), .ZN(n1844) );
  and2 U2048 ( .A1(n879), .A2(n1837), .Z(n1841) );
  inv1 U2049 ( .I(n879), .ZN(n1839) );
  and2 U2050 ( .A1(n1839), .A2(n1589), .Z(n1840) );
  or2 U2051 ( .A1(n1841), .A2(n1840), .Z(n1945) );
  inv1 U2052 ( .I(n1945), .ZN(n1842) );
  and2 U2053 ( .A1(f5), .A2(n1842), .Z(n1843) );
  or2 U2054 ( .A1(n1844), .A2(n1843), .Z(n1845) );
  and2 U2055 ( .A1(t5), .A2(n1845), .Z(n1846) );
  or2 U2056 ( .A1(n794), .A2(n1846), .Z(j10) );
  and2 U2057 ( .A1(a5), .A2(n189), .Z(n1847) );
  and2 U2058 ( .A1(n190), .A2(n1847), .Z(n1848) );
  or2 U2059 ( .A1(n1848), .A2(n109), .Z(n1874) );
  or2 U2061 ( .A1(n1850), .A2(n1880), .Z(n1858) );
  inv1 U2062 ( .I(n1850), .ZN(n1851) );
  or2 U2063 ( .A1(n1851), .A2(n1574), .Z(n1859) );
  or2 U2064 ( .A1(n1853), .A2(n1852), .Z(n1862) );
  or2 U2065 ( .A1(n1855), .A2(n1854), .Z(n1860) );
  and2 U2066 ( .A1(n1859), .A2(n1856), .Z(n1857) );
  and2 U2067 ( .A1(n1858), .A2(n1857), .Z(n1865) );
  and2 U2068 ( .A1(n1861), .A2(n1860), .Z(n1863) );
  and2 U2069 ( .A1(n1863), .A2(n1862), .Z(n1864) );
  or2 U2070 ( .A1(n1865), .A2(n1864), .Z(n1870) );
  and2 U2071 ( .A1(n726), .A2(n2019), .Z(n1868) );
  inv1 U2072 ( .I(n726), .ZN(n1866) );
  or2 U2074 ( .A1(n1868), .A2(n1867), .Z(n1881) );
  or2 U2076 ( .A1(n1870), .A2(n1879), .Z(n1869) );
  and2 U2077 ( .A1(n1874), .A2(n1869), .Z(n1873) );
  inv1 U2078 ( .I(n1870), .ZN(n1871) );
  or2 U2079 ( .A1(n1871), .A2(n1881), .Z(n1872) );
  inv1 U2081 ( .I(n1874), .ZN(n1892) );
  and2 U2082 ( .A1(n1876), .A2(n1875), .Z(n1878) );
  and2 U2083 ( .A1(n1113), .A2(n1571), .Z(n1877) );
  or2 U2084 ( .A1(n1878), .A2(n1877), .Z(n1895) );
  inv1 U2085 ( .I(n1895), .ZN(n1890) );
  and2 U2086 ( .A1(n1880), .A2(n1879), .Z(n1883) );
  and2 U2087 ( .A1(n1574), .A2(n1881), .Z(n1882) );
  or2 U2088 ( .A1(n1883), .A2(n1882), .Z(n1885) );
  and2 U2089 ( .A1(n1884), .A2(n1885), .Z(n1889) );
  and2 U2091 ( .A1(n1887), .A2(n1886), .Z(n1888) );
  or2 U2093 ( .A1(n1890), .A2(n1893), .Z(n1891) );
  and2 U2094 ( .A1(n1892), .A2(n1891), .Z(n1897) );
  inv1 U2095 ( .I(n1893), .ZN(n1894) );
  or2 U2096 ( .A1(n1895), .A2(n1894), .Z(n1896) );
  and2 U2097 ( .A1(n1897), .A2(n1896), .Z(n1898) );
  inv1 U2103 ( .I(n1917), .ZN(n1915) );
  inv1 U2104 ( .I(n644), .ZN(n1912) );
  and2 U2105 ( .A1(n645), .A2(n1912), .Z(n1906) );
  inv1 U2106 ( .I(n645), .ZN(n1904) );
  or2 U2108 ( .A1(n1906), .A2(n1905), .Z(n1907) );
  and2 U2109 ( .A1(n1915), .A2(n1907), .Z(n1910) );
  inv1 U2110 ( .I(n1907), .ZN(n1908) );
  and2 U2111 ( .A1(n1917), .A2(n1908), .Z(n1909) );
  and2 U2113 ( .A1(a5), .A2(n1928), .Z(n1922) );
  inv1 U2114 ( .I(n754), .ZN(n1911) );
  and2 U2115 ( .A1(n1911), .A2(n644), .Z(n1914) );
  and2 U2116 ( .A1(n754), .A2(n1912), .Z(n1913) );
  or2 U2117 ( .A1(n1914), .A2(n1913), .Z(n1916) );
  and2 U2118 ( .A1(n1916), .A2(n1915), .Z(n1920) );
  inv1 U2119 ( .I(n1916), .ZN(n1918) );
  and2 U2120 ( .A1(n1918), .A2(n1917), .Z(n1919) );
  and2 U2122 ( .A1(n1927), .A2(n1929), .Z(n1921) );
  or2 U2123 ( .A1(n1922), .A2(n1921), .Z(n1923) );
  and2 U2124 ( .A1(t5), .A2(n1923), .Z(n1924) );
  or2 U2125 ( .A1(n1924), .A2(n512), .Z(k10) );
  inv1 U2126 ( .I(u5), .ZN(n1926) );
  inv1 U2127 ( .I(l0), .ZN(n1925) );
  or2 U2128 ( .A1(n1926), .A2(n1925), .Z(n1937) );
  or2 U2129 ( .A1(n2022), .A2(n1939), .Z(n1935) );
  inv1 U2130 ( .I(a5), .ZN(n1927) );
  or2 U2134 ( .A1(n1933), .A2(n1932), .Z(n1934) );
  inv1 U2137 ( .I(n1970), .ZN(n1938) );
  and2 U2138 ( .A1(n1938), .A2(n53), .Z(n1950) );
  and2 U2139 ( .A1(k0), .A2(u5), .Z(n1942) );
  or2 U2140 ( .A1(n504), .A2(n1939), .Z(n1940) );
  inv1 U2141 ( .I(n1940), .ZN(n1941) );
  or2 U2142 ( .A1(n1942), .A2(n1941), .Z(n1948) );
  inv1 U2143 ( .I(f5), .ZN(n1944) );
  and2 U2145 ( .A1(f5), .A2(n1945), .Z(n1946) );
  and2 U2146 ( .A1(n1982), .A2(n1582), .Z(n1949) );
  or2 U2147 ( .A1(n1950), .A2(n1949), .Z(n1954) );
  and2 U2148 ( .A1(d), .A2(n1981), .Z(n1952) );
  and2 U2149 ( .A1(w), .A2(n52), .Z(n1951) );
  or2 U2150 ( .A1(n1952), .A2(n1951), .Z(n1953) );
  or2 U2151 ( .A1(n1954), .A2(n1953), .Z(l10) );
  and2 U2152 ( .A1(n15), .A2(w), .Z(n1956) );
  and2 U2153 ( .A1(n16), .A2(d), .Z(n1955) );
  or2 U2154 ( .A1(n1956), .A2(n1955), .Z(n1962) );
  and2 U2155 ( .A1(n1997), .A2(n1582), .Z(n1960) );
  or2 U2156 ( .A1(n1970), .A2(n1957), .Z(n1958) );
  inv1 U2157 ( .I(n1958), .ZN(n1959) );
  or2 U2158 ( .A1(n1960), .A2(n1959), .Z(n1961) );
  or2 U2159 ( .A1(n1962), .A2(n1961), .Z(m10) );
  or2 U2164 ( .A1(n2009), .A2(n408), .Z(n1966) );
  or2 U2165 ( .A1(n1966), .A2(n407), .Z(n1967) );
  inv1 U2167 ( .I(l1), .ZN(n1976) );
  or2 U2168 ( .A1(n1969), .A2(n1976), .Z(n10) );
  or2 U2169 ( .A1(n1583), .A2(d5), .Z(n1972) );
  or2 U2172 ( .A1(n2007), .A2(n322), .Z(n1974) );
  or2 U2173 ( .A1(n1974), .A2(n321), .Z(n1975) );
  inv1f U1654 ( .I(t3), .ZN(n1734) );
  inv1f U1655 ( .I(n1573), .ZN(n1574) );
  and2f U1656 ( .A1(x3), .A2(n1722), .Z(n1608) );
  or2f U1663 ( .A1(n1614), .A2(n1703), .Z(n1820) );
  or2 U1666 ( .A1(n1486), .A2(n1487), .Z(n661) );
  and2 U1669 ( .A1(n447), .A2(n1713), .Z(n1614) );
  inv1 U1670 ( .I(n648), .ZN(n647) );
  inv1 U1672 ( .I(n1901), .ZN(n1900) );
  and2f U1673 ( .A1(l2), .A2(n1734), .Z(n1686) );
  and2f U1680 ( .A1(c3), .A2(n1734), .Z(n1625) );
  and2f U1681 ( .A1(n2), .A2(n1734), .Z(n1653) );
  or2f U1688 ( .A1(n1808), .A2(n1779), .Z(n1663) );
  and2f U1689 ( .A1(p2), .A2(n1734), .Z(n1632) );
  inv1f U1691 ( .I(n729), .ZN(n1989) );
  or2f U1692 ( .A1(n1852), .A2(n1884), .Z(n729) );
  and2 U1693 ( .A1(n646), .A2(n647), .Z(n645) );
  inv1 U1702 ( .I(n1805), .ZN(n1804) );
  and2 U1728 ( .A1(n1866), .A2(n725), .Z(n1867) );
  inv1 U1729 ( .I(n1885), .ZN(n1886) );
  and2 U1732 ( .A1(n784), .A2(n691), .Z(n1486) );
  inv1 U1733 ( .I(n1887), .ZN(n1884) );
  or2 U1735 ( .A1(n1607), .A2(n1606), .Z(n1731) );
  inv1 U1738 ( .I(n1731), .ZN(n1729) );
  inv1 U1756 ( .I(n1838), .ZN(n1837) );
  and2 U1757 ( .A1(n1904), .A2(n644), .Z(n1905) );
  and2 U1774 ( .A1(n1991), .A2(n1901), .Z(n1902) );
  or2 U1778 ( .A1(n1666), .A2(n1665), .Z(n1794) );
  or2 U1801 ( .A1(n1568), .A2(n425), .Z(n1591) );
  or2 U1807 ( .A1(n1794), .A2(n425), .Z(n1753) );
  inv1f U1808 ( .I(s3), .ZN(n1722) );
  and2 U1809 ( .A1(m3), .A2(n1722), .Z(n1643) );
  and2f U1832 ( .A1(n1764), .A2(n1809), .Z(n1568) );
  or2 U1834 ( .A1(n1970), .A2(n2008), .Z(n1971) );
  or2f U1836 ( .A1(n1928), .A2(n1927), .Z(n1931) );
  inv1f U1838 ( .I(n1881), .ZN(n1879) );
  or2f U1839 ( .A1(n1818), .A2(n1819), .Z(n1838) );
  and2f U1849 ( .A1(n1944), .A2(n1943), .Z(n1947) );
  or2 U1854 ( .A1(n1583), .A2(b5), .Z(n1964) );
  and2f U1865 ( .A1(n669), .A2(n661), .Z(n1485) );
  or2f U1867 ( .A1(n1889), .A2(n1888), .Z(n1893) );
  inv1f U1868 ( .I(n1582), .ZN(n1583) );
  and2f U1869 ( .A1(n1833), .A2(n1832), .Z(n1834) );
  and2f U1895 ( .A1(n1793), .A2(n1792), .Z(n1819) );
  and2f U1924 ( .A1(n1788), .A2(n1787), .Z(n1793) );
  inv1f U1926 ( .I(n1764), .ZN(n1799) );
  or2f U2009 ( .A1(n1643), .A2(n1642), .Z(n1728) );
  inv1f U2012 ( .I(n1664), .ZN(n1666) );
  and2f U2015 ( .A1(n1931), .A2(n1930), .Z(n1933) );
  or2f U2017 ( .A1(n1929), .A2(a5), .Z(n1930) );
  or2f U2020 ( .A1(n1910), .A2(n1909), .Z(n1928) );
  and2f U2021 ( .A1(n678), .A2(n1900), .Z(n1903) );
  and2f U2026 ( .A1(n1572), .A2(n1689), .Z(n1571) );
  or2f U2028 ( .A1(n1574), .A2(n1887), .Z(n1689) );
  and2f U2029 ( .A1(n1972), .A2(n1971), .Z(n1973) );
  or2f U2030 ( .A1(n1899), .A2(n1898), .Z(n1901) );
  and2f U2031 ( .A1(n1873), .A2(n1872), .Z(n1899) );
  or2f U2032 ( .A1(n1819), .A2(n1818), .Z(n1589) );
  and2f U2035 ( .A1(n1964), .A2(n1963), .Z(n1965) );
  or2f U2037 ( .A1(n1970), .A2(n2010), .Z(n1963) );
  and2f U2040 ( .A1(n1797), .A2(n1593), .Z(n1592) );
  or2f U2042 ( .A1(n1796), .A2(n1809), .Z(n1797) );
  or2f U2044 ( .A1(n1829), .A2(n1828), .Z(n1833) );
  and2f U2045 ( .A1(n1825), .A2(n1824), .Z(n1829) );
  and2f U2060 ( .A1(n85), .A2(n1804), .Z(n1807) );
  and2f U2073 ( .A1(o3), .A2(n1722), .Z(n1606) );
  or2f U2075 ( .A1(n1729), .A2(n2014), .Z(n1780) );
  and2f U2080 ( .A1(n1968), .A2(n1967), .Z(n1969) );
  or2f U2090 ( .A1(n1965), .A2(c5), .Z(n1968) );
  or2f U2092 ( .A1(n1920), .A2(n1919), .Z(n1929) );
  or2f U2098 ( .A1(n1903), .A2(n1902), .Z(n1917) );
  and2f U2099 ( .A1(n1876), .A2(n1849), .Z(n1850) );
  and2f U2100 ( .A1(n1701), .A2(n1700), .Z(n1876) );
  or2f U2101 ( .A1(n1571), .A2(n1983), .Z(n1701) );
  and2f U2102 ( .A1(n1937), .A2(n1936), .Z(n1970) );
  and2f U2107 ( .A1(n1935), .A2(n1934), .Z(n1936) );
  or2f U2112 ( .A1(n1656), .A2(n1655), .Z(n1573) );
  or2f U2121 ( .A1(n1835), .A2(n1834), .Z(n1943) );
  and2f U2131 ( .A1(n1831), .A2(n1830), .Z(n1835) );
  or2f U2132 ( .A1(n1823), .A2(n1822), .Z(n1827) );
  and2f U2133 ( .A1(n1820), .A2(n1837), .Z(n1823) );
  and2f U2135 ( .A1(n425), .A2(n1588), .Z(n1803) );
  and2f U2136 ( .A1(n1797), .A2(n1593), .Z(n1588) );
  inv1f U2144 ( .I(n1668), .ZN(n1795) );
  or2f U2160 ( .A1(n1590), .A2(n1591), .Z(n1668) );
  and2f U2161 ( .A1(n1817), .A2(n1816), .Z(n1818) );
  and2f U2162 ( .A1(n1812), .A2(n1811), .Z(n1817) );
  or2f U2163 ( .A1(n1815), .A2(n1814), .Z(n1816) );
  and2f U2166 ( .A1(n1575), .A2(n1576), .Z(n1582) );
  or2f U2170 ( .A1(n1947), .A2(n1577), .Z(n1575) );
  or2f U2171 ( .A1(n1646), .A2(n1645), .Z(n1764) );
  and2f U2174 ( .A1(o4), .A2(n1730), .Z(n1646) );
endmodule

