
module b9 ( o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, 
        x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, 
        j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, 
        r0, q0, p0 );
  input o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w,
         v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0,
         s0, r0, q0, p0;
  wire   n186, n187, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n32, n33, n34, n38, n40, n43, n44, n49, n51, n66, n71,
         n73, n74, n75, n76, n77, n78, n85, n99, n102, n104, n105, n106, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n130, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n183, n184,
         n185, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197;

  and2 U13 ( .A1(l), .A2(n17), .Z(y0) );
  and2 U15 ( .A1(n18), .A2(d), .Z(w0) );
  and2 U16 ( .A1(n19), .A2(n20), .Z(n18) );
  or2 U17 ( .A1(n21), .A2(n22), .Z(n20) );
  and2 U19 ( .A1(z), .A2(n25), .Z(n24) );
  inv1 U20 ( .I(o), .ZN(n25) );
  and2 U21 ( .A1(a), .A2(n26), .Z(n23) );
  inv1 U22 ( .I(z), .ZN(n26) );
  inv1 U23 ( .I(m0), .ZN(n21) );
  inv1 U24 ( .I(n27), .ZN(n19) );
  and2 U25 ( .A1(n28), .A2(o), .Z(n27) );
  or2 U27 ( .A1(h0), .A2(f0), .Z(n30) );
  and2 U28 ( .A1(r), .A2(n183), .Z(n29) );
  inv1 U29 ( .I(n187), .ZN(v0) );
  or2 U30 ( .A1(n32), .A2(l0), .Z(n187) );
  and2 U31 ( .A1(c0), .A2(b0), .Z(n32) );
  or2 U32 ( .A1(v), .A2(n33), .Z(t0) );
  or2 U33 ( .A1(n33), .A2(n34), .Z(s0) );
  inv1 U34 ( .I(v), .ZN(n34) );
  inv1 U37 ( .I(l0), .ZN(n38) );
  inv1 U42 ( .I(n44), .ZN(n43) );
  or2 U43 ( .A1(c), .A2(d0), .Z(n44) );
  inv1 U48 ( .I(c), .ZN(n51) );
  inv1 U62 ( .I(i), .ZN(n49) );
  or2 U65 ( .A1(j), .A2(e0), .Z(n66) );
  and2 U70 ( .A1(b0), .A2(n190), .Z(n71) );
  and2 U75 ( .A1(n73), .A2(n74), .Z(g1) );
  and2 U76 ( .A1(b), .A2(n75), .Z(n74) );
  inv1 U77 ( .I(y), .ZN(n75) );
  and2 U78 ( .A1(x), .A2(w), .Z(n73) );
  and2 U79 ( .A1(n76), .A2(w), .Z(f1) );
  and2 U80 ( .A1(b), .A2(n77), .Z(n76) );
  inv1 U81 ( .I(x), .ZN(n77) );
  and2 U82 ( .A1(m), .A2(n17), .Z(e1) );
  and2 U83 ( .A1(n78), .A2(i0), .Z(n17) );
  and2 U84 ( .A1(a0), .A2(b0), .Z(n78) );
  or2 U91 ( .A1(t), .A2(s), .Z(n85) );
  or2 U121 ( .A1(n102), .A2(n192), .Z(p0) );
  inv1 U122 ( .I(n130), .ZN(n102) );
  or2 U124 ( .A1(n), .A2(e), .Z(n104) );
  and2 U125 ( .A1(n106), .A2(n195), .Z(n105) );
  inv1 U126 ( .I(n104), .ZN(n106) );
  inv1 U128 ( .I(n194), .ZN(n144) );
  buf0 U129 ( .I(n187), .Z(u0) );
  buf0 U130 ( .I(n195), .Z(x0) );
  buf0 U131 ( .I(n181), .Z(a1) );
  buf0 U132 ( .I(n185), .Z(c1) );
  buf0 U133 ( .I(n186), .Z(h1) );
  buf0 U134 ( .I(n181), .Z(i1) );
  inv1 U136 ( .I(j0), .ZN(n115) );
  and2 U137 ( .A1(c0), .A2(j0), .Z(n116) );
  or2 U138 ( .A1(n115), .A2(c0), .Z(n117) );
  inv1 U140 ( .I(e), .ZN(n184) );
  inv1 U141 ( .I(n116), .ZN(n119) );
  and2 U142 ( .A1(n119), .A2(b0), .Z(n122) );
  and2 U144 ( .A1(n188), .A2(n38), .Z(n121) );
  or2 U145 ( .A1(n122), .A2(n121), .Z(n33) );
  inv1 U146 ( .I(p), .ZN(n183) );
  inv1 U148 ( .I(n170), .ZN(n123) );
  or2 U149 ( .A1(n123), .A2(n189), .Z(n162) );
  and2 U153 ( .A1(k0), .A2(b0), .Z(n125) );
  or2 U154 ( .A1(n125), .A2(k), .Z(n126) );
  or2 U157 ( .A1(n144), .A2(e), .Z(n149) );
  or2 U158 ( .A1(n128), .A2(n114), .Z(n163) );
  inv1 U161 ( .I(n166), .ZN(n134) );
  inv1 U163 ( .I(k0), .ZN(n132) );
  and2 U166 ( .A1(n134), .A2(n142), .Z(n135) );
  or2 U167 ( .A1(n135), .A2(n184), .Z(q0) );
  and2 U168 ( .A1(e), .A2(n117), .Z(n136) );
  or2 U169 ( .A1(n136), .A2(n43), .Z(n141) );
  and2 U170 ( .A1(n188), .A2(e), .Z(n137) );
  or2 U171 ( .A1(n137), .A2(n51), .Z(n138) );
  and2 U172 ( .A1(n49), .A2(n138), .Z(n139) );
  or2 U173 ( .A1(n139), .A2(n144), .Z(n140) );
  or2 U174 ( .A1(n141), .A2(n140), .Z(r0) );
  and2 U177 ( .A1(n184), .A2(n196), .Z(n148) );
  and2 U178 ( .A1(f), .A2(n195), .Z(n146) );
  and2 U179 ( .A1(n144), .A2(h), .Z(n145) );
  or2 U180 ( .A1(n146), .A2(n145), .Z(n147) );
  inv1 U182 ( .I(n149), .ZN(n164) );
  and2 U183 ( .A1(f), .A2(n166), .Z(n150) );
  and2 U184 ( .A1(n164), .A2(n150), .Z(n153) );
  and2 U185 ( .A1(l0), .A2(b0), .Z(n151) );
  and2 U186 ( .A1(g), .A2(n151), .Z(n152) );
  or2 U187 ( .A1(n153), .A2(n152), .Z(n154) );
  inv1 U189 ( .I(n117), .ZN(n176) );
  and2 U190 ( .A1(i), .A2(n120), .Z(n157) );
  or2 U191 ( .A1(n157), .A2(n71), .Z(n158) );
  and2 U192 ( .A1(n176), .A2(n158), .Z(n161) );
  and2 U193 ( .A1(d0), .A2(i), .Z(n159) );
  and2 U194 ( .A1(n195), .A2(n159), .Z(n160) );
  inv1 U197 ( .I(n186), .ZN(n181) );
  and2 U198 ( .A1(n163), .A2(n162), .Z(b1) );
  inv1 U199 ( .I(c0), .ZN(n165) );
  or2 U202 ( .A1(n167), .A2(n99), .Z(n169) );
  and2 U203 ( .A1(n105), .A2(n169), .Z(n175) );
  and2 U204 ( .A1(u), .A2(b0), .Z(n173) );
  inv1 U205 ( .I(n85), .ZN(n171) );
  and2 U206 ( .A1(n171), .A2(n170), .Z(n172) );
  inv1 U209 ( .I(n185), .ZN(d1) );
  and2 U210 ( .A1(i), .A2(n176), .Z(n179) );
  or2 U212 ( .A1(n179), .A2(n178), .Z(n180) );
  inv1 U213 ( .I(n180), .ZN(j1) );
  inv1 U119 ( .I(n133), .ZN(n197) );
  and2 U120 ( .A1(n173), .A2(n172), .Z(n174) );
  inv1 U123 ( .I(n191), .ZN(n193) );
  inv1 U127 ( .I(n127), .ZN(n128) );
  and2 U135 ( .A1(n193), .A2(n127), .Z(n192) );
  inv1 U139 ( .I(b0), .ZN(n189) );
  inv1 U143 ( .I(b0), .ZN(n188) );
  inv1 U147 ( .I(b0), .ZN(n120) );
  or2f U150 ( .A1(n23), .A2(n24), .Z(n22) );
  or2f U151 ( .A1(n29), .A2(n30), .Z(n28) );
  inv1f U152 ( .I(e), .ZN(n190) );
  or2f U155 ( .A1(n175), .A2(n174), .Z(n185) );
  or2f U156 ( .A1(n155), .A2(n154), .Z(z0) );
  and2f U159 ( .A1(n148), .A2(n147), .Z(n155) );
  and2f U160 ( .A1(n165), .A2(b0), .Z(n168) );
  and2f U162 ( .A1(n124), .A2(q), .Z(n130) );
  or2f U164 ( .A1(n162), .A2(p), .Z(n124) );
  or2f U165 ( .A1(n161), .A2(n177), .Z(n186) );
  or2f U175 ( .A1(n160), .A2(n66), .Z(n177) );
  and2f U176 ( .A1(n156), .A2(n132), .Z(n133) );
  or2f U181 ( .A1(n115), .A2(c0), .Z(n156) );
  and2f U188 ( .A1(n118), .A2(k0), .Z(n167) );
  or2f U195 ( .A1(n118), .A2(n126), .Z(n127) );
  or2f U196 ( .A1(n177), .A2(n118), .Z(n178) );
  and2f U200 ( .A1(b0), .A2(j0), .Z(n118) );
  or2f U201 ( .A1(n168), .A2(n166), .Z(n99) );
  or2f U207 ( .A1(g0), .A2(e0), .Z(n166) );
  or2f U208 ( .A1(n40), .A2(l0), .Z(n170) );
  and2f U211 ( .A1(c0), .A2(j0), .Z(n40) );
  or2f U214 ( .A1(p), .A2(n114), .Z(n191) );
  or2f U215 ( .A1(n144), .A2(e), .Z(n114) );
  and2 U216 ( .A1(n0), .A2(o0), .Z(n195) );
  and2f U217 ( .A1(n0), .A2(o0), .Z(n194) );
  and2f U218 ( .A1(n197), .A2(b0), .Z(n196) );
  inv1 U219 ( .I(n196), .ZN(n142) );
endmodule

