
module C2670_iscas ( y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, 
        k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, 
        s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, 
        a6, z5, y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, 
        i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, 
        q4, p4, o4, n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, 
        y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, 
        g3, f3, e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, 
        o2, n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, 
        w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, 
        e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, 
        m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, 
        t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, i13, h13, 
        g13, f13, e13, d13, c13, b13, a13, z12, y12, x12, w12, v12, u12, t12, 
        s12, r12, q12, p12, o12, n12, m12, l12, k12, j12, i12, h12, g12, f12, 
        e12, d12, c12, b12, a12, z11, y11, x11, w11, v11, u11, t11, s11, r11, 
        q11, p11, o11, n11, m11, l11, k11, j11, i11, h11, g11, f11, e11, d11, 
        c11, b11, a11, z10, y10, x10, w10, v10, u10, t10, s10, r10, q10, p10, 
        o10, n10, m10, l10, k10, j10, i10, h10, g10, f10, e10, d10, c10, b10, 
        a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9, 
        j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8, s8, 
        r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8, b8, a8, 
        z7 );
  input y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, i7, h7,
         g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, q6,
         p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5,
         y5, x5, w5, v5, u5, t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5,
         h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4,
         q4, p4, o4, n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4,
         z3, y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3,
         i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2,
         r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, g2, f2, e2, d2, c2, b2,
         a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1,
         j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0,
         s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0,
         b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f,
         e, d, c, b, a;
  output i13, h13, g13, f13, e13, d13, c13, b13, a13, z12, y12, x12, w12, v12,
         u12, t12, s12, r12, q12, p12, o12, n12, m12, l12, k12, j12, i12, h12,
         g12, f12, e12, d12, c12, b12, a12, z11, y11, x11, w11, v11, u11, t11,
         s11, r11, q11, p11, o11, n11, m11, l11, k11, j11, i11, h11, g11, f11,
         e11, d11, c11, b11, a11, z10, y10, x10, w10, v10, u10, t10, s10, r10,
         q10, p10, o10, n10, m10, l10, k10, j10, i10, h10, g10, f10, e10, d10,
         c10, b10, a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9,
         l9, k9, j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8,
         u8, t8, s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8,
         d8, c8, b8, a8, z7;
  wire   e7, r6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5,
         t5, s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5,
         c5, b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4,
         l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3,
         u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, c281, f281, m281, a301,
         n9_snps_wire, n10_snps_wire, n12_snps_wire, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640;
  assign c11 = e7;
  assign d11 = e7;
  assign e11 = e7;
  assign a11 = r6;
  assign b11 = r6;
  assign x10 = i6;
  assign y10 = i6;
  assign z10 = i6;
  assign p11 = i6;
  assign w10 = h6;
  assign v10 = g6;
  assign u10 = f6;
  assign t10 = e6;
  assign s10 = d6;
  assign r10 = c6;
  assign q10 = b6;
  assign p10 = a6;
  assign o10 = z5;
  assign n10 = y5;
  assign m10 = x5;
  assign l10 = w5;
  assign k10 = v5;
  assign j10 = u5;
  assign i10 = t5;
  assign h10 = s5;
  assign g10 = r5;
  assign f10 = q5;
  assign e10 = p5;
  assign d10 = o5;
  assign c10 = n5;
  assign b10 = m5;
  assign a10 = l5;
  assign z9 = k5;
  assign y9 = j5;
  assign x9 = i5;
  assign w9 = h5;
  assign v9 = g5;
  assign u9 = f5;
  assign t9 = e5;
  assign s9 = d5;
  assign r9 = c5;
  assign q9 = b5;
  assign p9 = a5;
  assign o9 = z4;
  assign n9 = y4;
  assign m9 = x4;
  assign l9 = w4;
  assign k9 = v4;
  assign j9 = u4;
  assign i9 = t4;
  assign h9 = s4;
  assign g9 = r4;
  assign f9 = q4;
  assign e9 = p4;
  assign d9 = o4;
  assign c9 = n4;
  assign b9 = m4;
  assign a9 = l4;
  assign z8 = k4;
  assign y8 = j4;
  assign x8 = i4;
  assign w8 = h4;
  assign v8 = g4;
  assign u8 = f4;
  assign t8 = e4;
  assign s8 = d4;
  assign r8 = c4;
  assign q8 = b4;
  assign p8 = a4;
  assign o8 = z3;
  assign n8 = y3;
  assign m8 = x3;
  assign l8 = w3;
  assign k8 = v3;
  assign j8 = u3;
  assign i8 = t3;
  assign h8 = s3;
  assign g8 = r3;
  assign f8 = q3;
  assign e8 = p3;
  assign d8 = o3;
  assign c8 = n3;
  assign b8 = m3;
  assign a8 = l3;
  assign z7 = k3;
  assign n12 = c281;
  assign o12 = c281;
  assign p12 = f281;
  assign q12 = f281;
  assign s12 = m281;
  assign t12 = m281;
  assign c13 = a301;
  assign d13 = a301;
  assign g13 = 1'b0;

  inv1 U1 ( .I(y12), .ZN(z12) );
  and2 U2 ( .A1(n9_snps_wire), .A2(n10_snps_wire), .Z(y12) );
  and2 U3 ( .A1(n12_snps_wire), .A2(n13), .Z(n10_snps_wire) );
  or2 U4 ( .A1(w), .A2(n14), .Z(n13) );
  and2 U5 ( .A1(n15), .A2(n16), .Z(n14) );
  and2 U6 ( .A1(n17), .A2(n18), .Z(n16) );
  and2 U7 ( .A1(n19), .A2(n20), .Z(n18) );
  or2 U8 ( .A1(n21), .A2(n22), .Z(n20) );
  and2 U9 ( .A1(a0), .A2(n23), .Z(n22) );
  and2 U10 ( .A1(j7), .A2(n24), .Z(n21) );
  inv1 U11 ( .I(a0), .ZN(n24) );
  or2 U12 ( .A1(n25), .A2(n26), .Z(n19) );
  and2 U13 ( .A1(c7), .A2(n27), .Z(n26) );
  inv1 U14 ( .I(s), .ZN(n27) );
  and2 U15 ( .A1(s), .A2(n28), .Z(n25) );
  and2 U16 ( .A1(n29), .A2(n30), .Z(n17) );
  or2 U17 ( .A1(n31), .A2(n32), .Z(n30) );
  and2 U18 ( .A1(d7), .A2(n33), .Z(n32) );
  inv1 U19 ( .I(x), .ZN(n33) );
  and2 U20 ( .A1(x), .A2(n34), .Z(n31) );
  or2 U21 ( .A1(n35), .A2(n36), .Z(n29) );
  and2 U22 ( .A1(f7), .A2(n37), .Z(n36) );
  inv1 U23 ( .I(t), .ZN(n37) );
  and2 U24 ( .A1(t), .A2(n38), .Z(n35) );
  and2 U25 ( .A1(n39), .A2(n40), .Z(n15) );
  and2 U26 ( .A1(n41), .A2(n42), .Z(n40) );
  or2 U27 ( .A1(n43), .A2(n44), .Z(n42) );
  and2 U28 ( .A1(g7), .A2(n45), .Z(n44) );
  inv1 U29 ( .I(y), .ZN(n45) );
  and2 U30 ( .A1(y), .A2(n46), .Z(n43) );
  or2 U31 ( .A1(n47), .A2(n48), .Z(n41) );
  and2 U32 ( .A1(h7), .A2(n49), .Z(n48) );
  inv1 U33 ( .I(u), .ZN(n49) );
  and2 U34 ( .A1(u), .A2(n50), .Z(n47) );
  and2 U35 ( .A1(v), .A2(n51), .Z(n39) );
  or2 U36 ( .A1(n52), .A2(n53), .Z(n51) );
  and2 U37 ( .A1(i7), .A2(n54), .Z(n53) );
  inv1 U38 ( .I(z), .ZN(n54) );
  and2 U39 ( .A1(z), .A2(n55), .Z(n52) );
  and2 U40 ( .A1(n56), .A2(n57), .Z(n12_snps_wire) );
  or2 U41 ( .A1(l), .A2(n58), .Z(n57) );
  and2 U42 ( .A1(n59), .A2(n60), .Z(n58) );
  and2 U43 ( .A1(n61), .A2(n62), .Z(n60) );
  and2 U44 ( .A1(n63), .A2(n64), .Z(n62) );
  or2 U45 ( .A1(n65), .A2(n66), .Z(n64) );
  and2 U46 ( .A1(b7), .A2(n67), .Z(n66) );
  inv1 U47 ( .I(r), .ZN(n67) );
  and2 U48 ( .A1(r), .A2(n68), .Z(n65) );
  and2 U49 ( .A1(n69), .A2(n70), .Z(n63) );
  or2 U50 ( .A1(n71), .A2(n72), .Z(n70) );
  and2 U51 ( .A1(d), .A2(n73), .Z(n72) );
  and2 U52 ( .A1(t6), .A2(n74), .Z(n71) );
  inv1 U53 ( .I(d), .ZN(n74) );
  or2 U54 ( .A1(n75), .A2(n76), .Z(n69) );
  and2 U55 ( .A1(a7), .A2(n77), .Z(n76) );
  inv1 U56 ( .I(f), .ZN(n77) );
  and2 U57 ( .A1(f), .A2(n78), .Z(n75) );
  and2 U58 ( .A1(n79), .A2(n80), .Z(n61) );
  or2 U59 ( .A1(n81), .A2(n82), .Z(n80) );
  and2 U60 ( .A1(e), .A2(n83), .Z(n82) );
  and2 U61 ( .A1(w6), .A2(n84), .Z(n81) );
  inv1 U62 ( .I(e), .ZN(n84) );
  or2 U63 ( .A1(n85), .A2(n86), .Z(n79) );
  and2 U64 ( .A1(m), .A2(n87), .Z(n86) );
  and2 U65 ( .A1(s6), .A2(n88), .Z(n85) );
  inv1 U66 ( .I(m), .ZN(n88) );
  and2 U67 ( .A1(n89), .A2(n90), .Z(n59) );
  and2 U68 ( .A1(n91), .A2(n92), .Z(n90) );
  or2 U69 ( .A1(n93), .A2(n94), .Z(n92) );
  and2 U70 ( .A1(n), .A2(n95), .Z(n94) );
  and2 U71 ( .A1(v6), .A2(n96), .Z(n93) );
  inv1 U72 ( .I(n), .ZN(n96) );
  or2 U73 ( .A1(n97), .A2(n98), .Z(n91) );
  and2 U74 ( .A1(o), .A2(n99), .Z(n98) );
  and2 U75 ( .A1(x6), .A2(n100), .Z(n97) );
  inv1 U76 ( .I(o), .ZN(n100) );
  and2 U77 ( .A1(n101), .A2(n102), .Z(n89) );
  or2 U78 ( .A1(n103), .A2(n104), .Z(n102) );
  and2 U79 ( .A1(p), .A2(n105), .Z(n104) );
  and2 U80 ( .A1(y6), .A2(n106), .Z(n103) );
  inv1 U81 ( .I(p), .ZN(n106) );
  or2 U82 ( .A1(n107), .A2(n108), .Z(n101) );
  and2 U83 ( .A1(q), .A2(n109), .Z(n108) );
  and2 U84 ( .A1(z6), .A2(n110), .Z(n107) );
  inv1 U85 ( .I(q), .ZN(n110) );
  or2 U86 ( .A1(n111), .A2(n112), .Z(n56) );
  inv1 U87 ( .I(l), .ZN(n112) );
  and2 U88 ( .A1(n113), .A2(n114), .Z(n111) );
  and2 U89 ( .A1(n115), .A2(n116), .Z(n114) );
  and2 U90 ( .A1(n117), .A2(n118), .Z(n116) );
  and2 U91 ( .A1(n119), .A2(n120), .Z(n118) );
  or2 U92 ( .A1(n121), .A2(n73), .Z(n120) );
  or2 U93 ( .A1(t6), .A2(n122), .Z(n119) );
  and2 U94 ( .A1(n123), .A2(n124), .Z(n117) );
  and2 U95 ( .A1(n125), .A2(n126), .Z(n124) );
  or2 U96 ( .A1(n127), .A2(n95), .Z(n126) );
  or2 U97 ( .A1(v6), .A2(g12), .Z(n125) );
  and2 U98 ( .A1(n128), .A2(n129), .Z(n123) );
  or2 U99 ( .A1(n130), .A2(n87), .Z(n129) );
  or2 U100 ( .A1(s6), .A2(n131), .Z(n128) );
  and2 U101 ( .A1(n132), .A2(n133), .Z(n115) );
  and2 U102 ( .A1(n134), .A2(n135), .Z(n133) );
  or2 U103 ( .A1(c12), .A2(n83), .Z(n135) );
  or2 U104 ( .A1(w6), .A2(h12), .Z(n134) );
  and2 U105 ( .A1(n136), .A2(n137), .Z(n132) );
  or2 U106 ( .A1(b12), .A2(n99), .Z(n137) );
  or2 U107 ( .A1(x6), .A2(i12), .Z(n136) );
  and2 U108 ( .A1(n138), .A2(n139), .Z(n113) );
  and2 U109 ( .A1(n140), .A2(n141), .Z(n139) );
  and2 U110 ( .A1(n142), .A2(n143), .Z(n141) );
  or2 U111 ( .A1(a12), .A2(n105), .Z(n143) );
  or2 U112 ( .A1(y6), .A2(j12), .Z(n142) );
  and2 U113 ( .A1(n144), .A2(n145), .Z(n140) );
  or2 U114 ( .A1(n146), .A2(n109), .Z(n145) );
  or2 U115 ( .A1(z6), .A2(k12), .Z(n144) );
  and2 U116 ( .A1(n147), .A2(n148), .Z(n138) );
  and2 U117 ( .A1(n149), .A2(n150), .Z(n148) );
  or2 U118 ( .A1(n151), .A2(n78), .Z(n150) );
  or2 U119 ( .A1(a7), .A2(l12), .Z(n149) );
  and2 U120 ( .A1(n152), .A2(n153), .Z(n147) );
  or2 U121 ( .A1(n154), .A2(n68), .Z(n153) );
  or2 U122 ( .A1(b7), .A2(m12), .Z(n152) );
  and2 U123 ( .A1(i), .A2(n155), .Z(n9_snps_wire) );
  or2 U124 ( .A1(n156), .A2(n157), .Z(n155) );
  inv1 U125 ( .I(w), .ZN(n157) );
  and2 U126 ( .A1(n158), .A2(n159), .Z(n156) );
  and2 U127 ( .A1(n160), .A2(n161), .Z(n159) );
  and2 U128 ( .A1(n162), .A2(n163), .Z(n161) );
  and2 U129 ( .A1(n164), .A2(n165), .Z(n162) );
  or2 U130 ( .A1(y11), .A2(n23), .Z(n165) );
  or2 U131 ( .A1(j7), .A2(n166), .Z(n164) );
  and2 U132 ( .A1(n167), .A2(n168), .Z(n160) );
  and2 U133 ( .A1(n169), .A2(n170), .Z(n168) );
  or2 U134 ( .A1(x11), .A2(n55), .Z(n170) );
  or2 U135 ( .A1(i7), .A2(n171), .Z(n169) );
  and2 U136 ( .A1(n172), .A2(n173), .Z(n167) );
  or2 U137 ( .A1(z11), .A2(n50), .Z(n173) );
  or2 U138 ( .A1(h7), .A2(n174), .Z(n172) );
  and2 U139 ( .A1(n175), .A2(n176), .Z(n158) );
  and2 U140 ( .A1(n177), .A2(n178), .Z(n176) );
  and2 U141 ( .A1(n179), .A2(n180), .Z(n178) );
  or2 U142 ( .A1(n181), .A2(n46), .Z(n180) );
  or2 U143 ( .A1(g7), .A2(n182), .Z(n179) );
  and2 U144 ( .A1(n183), .A2(n184), .Z(n177) );
  or2 U145 ( .A1(n185), .A2(n28), .Z(n184) );
  or2 U146 ( .A1(c7), .A2(n186), .Z(n183) );
  and2 U147 ( .A1(n187), .A2(n188), .Z(n175) );
  and2 U148 ( .A1(n189), .A2(n190), .Z(n188) );
  or2 U149 ( .A1(n191), .A2(n38), .Z(n190) );
  or2 U150 ( .A1(f7), .A2(n192), .Z(n189) );
  and2 U151 ( .A1(n193), .A2(n194), .Z(n187) );
  or2 U152 ( .A1(n195), .A2(n34), .Z(n194) );
  or2 U153 ( .A1(d7), .A2(n196), .Z(n193) );
  or2 U154 ( .A1(l7), .A2(n197), .Z(u12) );
  or2 U155 ( .A1(n198), .A2(n199), .Z(n197) );
  and2 U156 ( .A1(n200), .A2(n201), .Z(n199) );
  and2 U157 ( .A1(k7), .A2(n163), .Z(n198) );
  inv1 U158 ( .I(v11), .ZN(u11) );
  or2 U159 ( .A1(n202), .A2(n203), .Z(v11) );
  or2 U160 ( .A1(r11), .A2(n204), .Z(t11) );
  inv1 U161 ( .I(o7), .ZN(n204) );
  or2 U162 ( .A1(r11), .A2(n205), .Z(s11) );
  inv1 U163 ( .I(m6), .ZN(n205) );
  or2 U164 ( .A1(n206), .A2(n122), .Z(r12) );
  and2 U165 ( .A1(n207), .A2(n208), .Z(n206) );
  inv1 U166 ( .I(n209), .ZN(r11) );
  and2 U167 ( .A1(g), .A2(o6), .Z(n209) );
  and2 U168 ( .A1(v1), .A2(i6), .Z(q11) );
  inv1 U169 ( .I(n210), .ZN(o11) );
  and2 U170 ( .A1(n211), .A2(k), .Z(n210) );
  and2 U171 ( .A1(b), .A2(o6), .Z(n211) );
  or2 U172 ( .A1(n212), .A2(n213), .Z(n11) );
  or2 U173 ( .A1(n50), .A2(n55), .Z(n213) );
  or2 U174 ( .A1(n23), .A2(n46), .Z(n212) );
  or2 U175 ( .A1(n214), .A2(n215), .Z(m281) );
  and2 U176 ( .A1(n131), .A2(n216), .Z(n215) );
  and2 U177 ( .A1(q6), .A2(n207), .Z(n214) );
  inv1 U178 ( .I(i13), .ZN(h13) );
  or2 U179 ( .A1(n217), .A2(n218), .Z(i13) );
  or2 U180 ( .A1(n219), .A2(n220), .Z(n218) );
  or2 U181 ( .A1(x12), .A2(w12), .Z(n220) );
  and2 U182 ( .A1(n221), .A2(n222), .Z(w12) );
  inv1 U183 ( .I(n223), .ZN(n222) );
  and2 U184 ( .A1(n224), .A2(n225), .Z(n223) );
  or2 U185 ( .A1(n225), .A2(n224), .Z(n221) );
  or2 U186 ( .A1(n226), .A2(n227), .Z(n224) );
  inv1 U187 ( .I(n228), .ZN(n227) );
  or2 U188 ( .A1(n229), .A2(n230), .Z(n228) );
  and2 U189 ( .A1(n230), .A2(n229), .Z(n226) );
  inv1 U190 ( .I(n231), .ZN(n229) );
  or2 U191 ( .A1(n232), .A2(n233), .Z(n231) );
  and2 U192 ( .A1(f7), .A2(n46), .Z(n233) );
  and2 U193 ( .A1(g7), .A2(n38), .Z(n232) );
  or2 U194 ( .A1(n234), .A2(n235), .Z(n230) );
  and2 U195 ( .A1(h7), .A2(n55), .Z(n235) );
  inv1 U196 ( .I(i7), .ZN(n55) );
  and2 U197 ( .A1(i7), .A2(n50), .Z(n234) );
  and2 U198 ( .A1(n236), .A2(n237), .Z(n225) );
  inv1 U199 ( .I(n238), .ZN(n237) );
  and2 U200 ( .A1(n239), .A2(n240), .Z(n238) );
  or2 U201 ( .A1(n240), .A2(n239), .Z(n236) );
  or2 U202 ( .A1(n241), .A2(n242), .Z(n239) );
  and2 U203 ( .A1(j7), .A2(n201), .Z(n242) );
  inv1 U204 ( .I(k7), .ZN(n201) );
  and2 U205 ( .A1(k7), .A2(n23), .Z(n241) );
  inv1 U206 ( .I(j7), .ZN(n23) );
  and2 U207 ( .A1(n243), .A2(n244), .Z(n240) );
  or2 U208 ( .A1(n245), .A2(y7), .Z(n244) );
  inv1 U209 ( .I(n246), .ZN(n243) );
  and2 U210 ( .A1(y7), .A2(n245), .Z(n246) );
  inv1 U211 ( .I(l7), .ZN(n245) );
  and2 U212 ( .A1(n247), .A2(n248), .Z(x12) );
  or2 U213 ( .A1(n249), .A2(n250), .Z(n248) );
  inv1 U214 ( .I(n251), .ZN(n247) );
  and2 U215 ( .A1(n250), .A2(n249), .Z(n251) );
  and2 U216 ( .A1(n252), .A2(n253), .Z(n249) );
  or2 U217 ( .A1(n254), .A2(b7), .Z(n253) );
  or2 U218 ( .A1(n68), .A2(n255), .Z(n252) );
  inv1 U219 ( .I(n254), .ZN(n255) );
  and2 U220 ( .A1(n256), .A2(n257), .Z(n254) );
  or2 U221 ( .A1(n258), .A2(n259), .Z(n257) );
  inv1 U222 ( .I(n260), .ZN(n259) );
  or2 U223 ( .A1(n260), .A2(n261), .Z(n256) );
  inv1 U224 ( .I(n258), .ZN(n261) );
  and2 U225 ( .A1(n262), .A2(n263), .Z(n258) );
  or2 U226 ( .A1(n264), .A2(a7), .Z(n263) );
  inv1 U227 ( .I(n265), .ZN(n264) );
  or2 U228 ( .A1(n78), .A2(n265), .Z(n262) );
  or2 U229 ( .A1(n266), .A2(n267), .Z(n265) );
  and2 U230 ( .A1(v6), .A2(n83), .Z(n267) );
  and2 U231 ( .A1(w6), .A2(n95), .Z(n266) );
  and2 U232 ( .A1(n268), .A2(n269), .Z(n260) );
  or2 U233 ( .A1(n270), .A2(n271), .Z(n269) );
  inv1 U234 ( .I(n272), .ZN(n268) );
  and2 U235 ( .A1(n271), .A2(n270), .Z(n272) );
  and2 U236 ( .A1(n273), .A2(n274), .Z(n270) );
  or2 U237 ( .A1(n99), .A2(x7), .Z(n274) );
  inv1 U238 ( .I(x6), .ZN(n99) );
  or2 U239 ( .A1(n275), .A2(x6), .Z(n273) );
  inv1 U240 ( .I(x7), .ZN(n275) );
  or2 U241 ( .A1(n276), .A2(n277), .Z(n271) );
  and2 U242 ( .A1(y6), .A2(n109), .Z(n277) );
  and2 U243 ( .A1(z6), .A2(n105), .Z(n276) );
  inv1 U244 ( .I(y6), .ZN(n105) );
  or2 U245 ( .A1(n278), .A2(n279), .Z(n250) );
  and2 U246 ( .A1(c7), .A2(n34), .Z(n279) );
  and2 U247 ( .A1(d7), .A2(n28), .Z(n278) );
  or2 U248 ( .A1(e13), .A2(n280), .Z(n217) );
  or2 U249 ( .A1(v12), .A2(b13), .Z(n280) );
  and2 U250 ( .A1(j), .A2(n281), .Z(v12) );
  and2 U251 ( .A1(n282), .A2(n283), .Z(n281) );
  or2 U252 ( .A1(n284), .A2(n285), .Z(n283) );
  inv1 U253 ( .I(n286), .ZN(n282) );
  and2 U254 ( .A1(n285), .A2(n284), .Z(n286) );
  and2 U255 ( .A1(n287), .A2(n288), .Z(n284) );
  or2 U256 ( .A1(n289), .A2(t6), .Z(n288) );
  or2 U257 ( .A1(n73), .A2(n290), .Z(n287) );
  inv1 U258 ( .I(n289), .ZN(n290) );
  and2 U259 ( .A1(n291), .A2(n292), .Z(n289) );
  inv1 U260 ( .I(n293), .ZN(n292) );
  and2 U261 ( .A1(n294), .A2(n295), .Z(n293) );
  or2 U262 ( .A1(n295), .A2(n294), .Z(n291) );
  or2 U263 ( .A1(n296), .A2(n297), .Z(n294) );
  inv1 U264 ( .I(n298), .ZN(n297) );
  or2 U265 ( .A1(n299), .A2(p7), .Z(n298) );
  and2 U266 ( .A1(p7), .A2(n299), .Z(n296) );
  and2 U267 ( .A1(n300), .A2(n301), .Z(n299) );
  or2 U268 ( .A1(n302), .A2(r7), .Z(n301) );
  inv1 U269 ( .I(n303), .ZN(n300) );
  and2 U270 ( .A1(r7), .A2(n302), .Z(n303) );
  inv1 U271 ( .I(q7), .ZN(n302) );
  and2 U272 ( .A1(n304), .A2(n305), .Z(n295) );
  inv1 U273 ( .I(n306), .ZN(n305) );
  and2 U274 ( .A1(n307), .A2(n308), .Z(n306) );
  or2 U275 ( .A1(n308), .A2(n307), .Z(n304) );
  or2 U276 ( .A1(n309), .A2(n310), .Z(n307) );
  and2 U277 ( .A1(s6), .A2(n311), .Z(n310) );
  inv1 U278 ( .I(s7), .ZN(n311) );
  and2 U279 ( .A1(s7), .A2(n87), .Z(n309) );
  and2 U280 ( .A1(n312), .A2(n313), .Z(n308) );
  or2 U281 ( .A1(n314), .A2(u7), .Z(n313) );
  inv1 U282 ( .I(t7), .ZN(n314) );
  or2 U283 ( .A1(n315), .A2(t7), .Z(n312) );
  inv1 U284 ( .I(u7), .ZN(n315) );
  or2 U285 ( .A1(n316), .A2(n317), .Z(n285) );
  inv1 U286 ( .I(n318), .ZN(n317) );
  or2 U287 ( .A1(n319), .A2(w7), .Z(n318) );
  and2 U288 ( .A1(w7), .A2(n319), .Z(n316) );
  inv1 U289 ( .I(v7), .ZN(n319) );
  or2 U291 ( .A1(n320), .A2(n321), .Z(f281) );
  and2 U292 ( .A1(q6), .A2(i12), .Z(n321) );
  and2 U293 ( .A1(g12), .A2(n216), .Z(n320) );
  and2 U295 ( .A1(n324), .A2(n325), .Z(n323) );
  and2 U298 ( .A1(n330), .A2(n331), .Z(n329) );
  or2 U301 ( .A1(n336), .A2(n337), .Z(n335) );
  and2 U302 ( .A1(n338), .A2(n339), .Z(n337) );
  and2 U303 ( .A1(n340), .A2(n341), .Z(n338) );
  or2 U305 ( .A1(n343), .A2(n344), .Z(n340) );
  and2 U308 ( .A1(n349), .A2(n350), .Z(n348) );
  and2 U311 ( .A1(n355), .A2(n356), .Z(n354) );
  and2 U314 ( .A1(n361), .A2(n362), .Z(n360) );
  and2 U317 ( .A1(n367), .A2(n368), .Z(n366) );
  and2 U320 ( .A1(n373), .A2(n374), .Z(n372) );
  or2 U323 ( .A1(n376), .A2(n377), .Z(n374) );
  and2 U324 ( .A1(n378), .A2(n83), .Z(n377) );
  inv1 U325 ( .I(w6), .ZN(n83) );
  and2 U326 ( .A1(n379), .A2(n50), .Z(n376) );
  inv1 U327 ( .I(h7), .ZN(n50) );
  and2 U329 ( .A1(n382), .A2(n127), .Z(n381) );
  or2 U331 ( .A1(n385), .A2(n386), .Z(n384) );
  and2 U332 ( .A1(n387), .A2(n121), .Z(n386) );
  and2 U333 ( .A1(n388), .A2(n130), .Z(n385) );
  and2 U334 ( .A1(n389), .A2(n390), .Z(n388) );
  or2 U335 ( .A1(n391), .A2(n392), .Z(n390) );
  inv1 U337 ( .I(s6), .ZN(n87) );
  or2 U339 ( .A1(n121), .A2(n387), .Z(n389) );
  inv1 U342 ( .I(t6), .ZN(n73) );
  or2 U344 ( .A1(n127), .A2(n382), .Z(n383) );
  or2 U345 ( .A1(n395), .A2(n396), .Z(n382) );
  and2 U346 ( .A1(n378), .A2(n95), .Z(n396) );
  inv1 U347 ( .I(v6), .ZN(n95) );
  and2 U348 ( .A1(n379), .A2(n46), .Z(n395) );
  inv1 U349 ( .I(g7), .ZN(n46) );
  or2 U350 ( .A1(n367), .A2(n368), .Z(n369) );
  or2 U351 ( .A1(b12), .A2(n397), .Z(n368) );
  inv1 U352 ( .I(n398), .ZN(n367) );
  or2 U353 ( .A1(n397), .A2(n399), .Z(n398) );
  or2 U354 ( .A1(n400), .A2(n401), .Z(n399) );
  and2 U355 ( .A1(x6), .A2(n378), .Z(n401) );
  and2 U356 ( .A1(n379), .A2(i7), .Z(n400) );
  or2 U357 ( .A1(n361), .A2(n362), .Z(n363) );
  or2 U358 ( .A1(a12), .A2(n397), .Z(n362) );
  inv1 U359 ( .I(n402), .ZN(n361) );
  or2 U360 ( .A1(n397), .A2(n403), .Z(n402) );
  or2 U361 ( .A1(n404), .A2(n405), .Z(n403) );
  and2 U362 ( .A1(y6), .A2(n378), .Z(n405) );
  and2 U363 ( .A1(n379), .A2(j7), .Z(n404) );
  inv1 U364 ( .I(h), .ZN(n397) );
  or2 U365 ( .A1(n355), .A2(n356), .Z(n357) );
  or2 U366 ( .A1(n146), .A2(n406), .Z(n356) );
  and2 U367 ( .A1(n109), .A2(n407), .Z(n355) );
  inv1 U368 ( .I(z6), .ZN(n109) );
  or2 U369 ( .A1(n349), .A2(n350), .Z(n351) );
  or2 U370 ( .A1(n151), .A2(n406), .Z(n350) );
  inv1 U371 ( .I(n407), .ZN(n406) );
  and2 U372 ( .A1(n78), .A2(n407), .Z(n349) );
  and2 U373 ( .A1(n378), .A2(h), .Z(n407) );
  inv1 U378 ( .I(u6), .ZN(n410) );
  inv1 U379 ( .I(a7), .ZN(n78) );
  or2 U380 ( .A1(n339), .A2(n341), .Z(n345) );
  or2 U381 ( .A1(n154), .A2(n411), .Z(n341) );
  and2 U382 ( .A1(n68), .A2(n412), .Z(n339) );
  inv1 U383 ( .I(b7), .ZN(n68) );
  and2 U384 ( .A1(n343), .A2(n344), .Z(n334) );
  or2 U385 ( .A1(n185), .A2(n411), .Z(n344) );
  and2 U386 ( .A1(n28), .A2(n412), .Z(n343) );
  inv1 U387 ( .I(c7), .ZN(n28) );
  or2 U388 ( .A1(n330), .A2(n331), .Z(n332) );
  or2 U389 ( .A1(n195), .A2(n411), .Z(n331) );
  and2 U390 ( .A1(n34), .A2(n412), .Z(n330) );
  inv1 U391 ( .I(d7), .ZN(n34) );
  or2 U392 ( .A1(n324), .A2(n325), .Z(n326) );
  or2 U393 ( .A1(n191), .A2(n411), .Z(n325) );
  inv1 U394 ( .I(n412), .ZN(n411) );
  and2 U395 ( .A1(n38), .A2(n412), .Z(n324) );
  and2 U396 ( .A1(d0), .A2(n413), .Z(n412) );
  and2 U397 ( .A1(n414), .A2(x11), .Z(n413) );
  or2 U398 ( .A1(z11), .A2(u6), .Z(n414) );
  inv1 U399 ( .I(f7), .ZN(n38) );
  or2 U400 ( .A1(n415), .A2(n416), .Z(f12) );
  and2 U401 ( .A1(c), .A2(a), .Z(n415) );
  inv1 U402 ( .I(n417), .ZN(e13) );
  or2 U403 ( .A1(c0), .A2(n418), .Z(n417) );
  or2 U404 ( .A1(n419), .A2(n420), .Z(n418) );
  inv1 U405 ( .I(n421), .ZN(n420) );
  or2 U406 ( .A1(n422), .A2(n423), .Z(n421) );
  and2 U407 ( .A1(n423), .A2(n422), .Z(n419) );
  and2 U408 ( .A1(n424), .A2(n425), .Z(n422) );
  or2 U409 ( .A1(n426), .A2(n427), .Z(n425) );
  inv1 U410 ( .I(n428), .ZN(n424) );
  and2 U411 ( .A1(n427), .A2(n426), .Z(n428) );
  or2 U412 ( .A1(n429), .A2(n430), .Z(n423) );
  and2 U413 ( .A1(i12), .A2(c12), .Z(n430) );
  and2 U414 ( .A1(h12), .A2(b12), .Z(n429) );
  or2 U415 ( .A1(n416), .A2(n431), .Z(e12) );
  inv1 U416 ( .I(b0), .ZN(n431) );
  inv1 U417 ( .I(n432), .ZN(n416) );
  and2 U418 ( .A1(j6), .A2(n433), .Z(n432) );
  and2 U419 ( .A1(o6), .A2(w11), .Z(n433) );
  inv1 U420 ( .I(n219), .ZN(w11) );
  or2 U421 ( .A1(n434), .A2(n435), .Z(n219) );
  and2 U422 ( .A1(m6), .A2(n202), .Z(n435) );
  or2 U423 ( .A1(n436), .A2(n437), .Z(n202) );
  or2 U424 ( .A1(k11), .A2(j11), .Z(n437) );
  inv1 U425 ( .I(a1), .ZN(j11) );
  inv1 U426 ( .I(r2), .ZN(k11) );
  or2 U427 ( .A1(m11), .A2(l11), .Z(n436) );
  inv1 U428 ( .I(q0), .ZN(l11) );
  inv1 U429 ( .I(h2), .ZN(m11) );
  and2 U430 ( .A1(o7), .A2(n203), .Z(n434) );
  or2 U431 ( .A1(n438), .A2(n439), .Z(n203) );
  or2 U432 ( .A1(g11), .A2(f11), .Z(n439) );
  inv1 U433 ( .I(f0), .ZN(f11) );
  inv1 U434 ( .I(b3), .ZN(g11) );
  or2 U435 ( .A1(i11), .A2(h11), .Z(n438) );
  inv1 U436 ( .I(l1), .ZN(h11) );
  inv1 U437 ( .I(x1), .ZN(i11) );
  or2 U438 ( .A1(n131), .A2(n208), .Z(d12) );
  inv1 U439 ( .I(p6), .ZN(n208) );
  or2 U440 ( .A1(n440), .A2(n441), .Z(c281) );
  and2 U441 ( .A1(q6), .A2(h12), .Z(n441) );
  and2 U442 ( .A1(n122), .A2(n216), .Z(n440) );
  inv1 U443 ( .I(h12), .ZN(c12) );
  or2 U444 ( .A1(n442), .A2(n443), .Z(h12) );
  or2 U445 ( .A1(n444), .A2(n445), .Z(n443) );
  and2 U446 ( .A1(v0), .A2(n446), .Z(n445) );
  and2 U447 ( .A1(l0), .A2(n447), .Z(n444) );
  or2 U448 ( .A1(n448), .A2(n449), .Z(n442) );
  and2 U449 ( .A1(g1), .A2(n450), .Z(n449) );
  and2 U450 ( .A1(r1), .A2(n451), .Z(n448) );
  inv1 U451 ( .I(n452), .ZN(b13) );
  or2 U452 ( .A1(c0), .A2(n453), .Z(n452) );
  or2 U453 ( .A1(n454), .A2(n455), .Z(n453) );
  and2 U454 ( .A1(n456), .A2(n457), .Z(n455) );
  inv1 U455 ( .I(n458), .ZN(n454) );
  or2 U456 ( .A1(n457), .A2(n456), .Z(n458) );
  or2 U457 ( .A1(n459), .A2(n460), .Z(n456) );
  and2 U458 ( .A1(x11), .A2(n163), .Z(n460) );
  and2 U460 ( .A1(n200), .A2(n171), .Z(n459) );
  inv1 U468 ( .I(n163), .ZN(n200) );
  or2 U469 ( .A1(n471), .A2(n472), .Z(n163) );
  or2 U470 ( .A1(n473), .A2(n474), .Z(n472) );
  and2 U471 ( .A1(i2), .A2(n465), .Z(n474) );
  and2 U472 ( .A1(s2), .A2(n466), .Z(n473) );
  or2 U473 ( .A1(n475), .A2(n476), .Z(n471) );
  and2 U474 ( .A1(y1), .A2(n469), .Z(n476) );
  and2 U475 ( .A1(c3), .A2(n470), .Z(n475) );
  and2 U476 ( .A1(n477), .A2(n478), .Z(n457) );
  inv1 U477 ( .I(n479), .ZN(n478) );
  and2 U478 ( .A1(n480), .A2(n481), .Z(n479) );
  or2 U479 ( .A1(n481), .A2(n480), .Z(n477) );
  or2 U480 ( .A1(n482), .A2(n483), .Z(n480) );
  and2 U481 ( .A1(n484), .A2(n485), .Z(n483) );
  inv1 U482 ( .I(n486), .ZN(n482) );
  or2 U483 ( .A1(n485), .A2(n484), .Z(n486) );
  or2 U484 ( .A1(n487), .A2(n488), .Z(n484) );
  and2 U485 ( .A1(y11), .A2(n174), .Z(n488) );
  inv1 U486 ( .I(n166), .ZN(y11) );
  and2 U487 ( .A1(z11), .A2(n166), .Z(n487) );
  or2 U488 ( .A1(n489), .A2(n490), .Z(n166) );
  or2 U489 ( .A1(n491), .A2(n492), .Z(n490) );
  and2 U490 ( .A1(j2), .A2(n465), .Z(n492) );
  and2 U491 ( .A1(t2), .A2(n466), .Z(n491) );
  or2 U492 ( .A1(n493), .A2(n494), .Z(n489) );
  and2 U493 ( .A1(z1), .A2(n469), .Z(n494) );
  and2 U494 ( .A1(d3), .A2(n470), .Z(n493) );
  inv1 U495 ( .I(n174), .ZN(z11) );
  or2 U497 ( .A1(n497), .A2(n498), .Z(n496) );
  or2 U503 ( .A1(n501), .A2(n502), .Z(n485) );
  or2 U504 ( .A1(n503), .A2(n504), .Z(n502) );
  and2 U505 ( .A1(p2), .A2(n465), .Z(n504) );
  and2 U506 ( .A1(z2), .A2(n466), .Z(n503) );
  or2 U507 ( .A1(n505), .A2(n506), .Z(n501) );
  and2 U508 ( .A1(f2), .A2(n469), .Z(n506) );
  and2 U509 ( .A1(j3), .A2(n470), .Z(n505) );
  and2 U510 ( .A1(n507), .A2(n508), .Z(n481) );
  or2 U511 ( .A1(n509), .A2(n510), .Z(n508) );
  inv1 U512 ( .I(n511), .ZN(n507) );
  and2 U513 ( .A1(n510), .A2(n509), .Z(n511) );
  inv1 U514 ( .I(n512), .ZN(n509) );
  or2 U515 ( .A1(n513), .A2(n514), .Z(n512) );
  and2 U516 ( .A1(n181), .A2(n186), .Z(n514) );
  inv1 U517 ( .I(n182), .ZN(n181) );
  and2 U518 ( .A1(n185), .A2(n182), .Z(n513) );
  or2 U519 ( .A1(n515), .A2(n516), .Z(n182) );
  or2 U520 ( .A1(n517), .A2(n518), .Z(n516) );
  and2 U521 ( .A1(m2), .A2(n465), .Z(n518) );
  and2 U522 ( .A1(w2), .A2(n466), .Z(n517) );
  or2 U523 ( .A1(n519), .A2(n520), .Z(n515) );
  and2 U524 ( .A1(c2), .A2(n469), .Z(n520) );
  and2 U525 ( .A1(g3), .A2(n470), .Z(n519) );
  inv1 U526 ( .I(n186), .ZN(n185) );
  or2 U527 ( .A1(n521), .A2(n522), .Z(n186) );
  or2 U528 ( .A1(n523), .A2(n524), .Z(n522) );
  and2 U529 ( .A1(g2), .A2(n465), .Z(n524) );
  and2 U530 ( .A1(q2), .A2(n466), .Z(n523) );
  or2 U531 ( .A1(n525), .A2(n526), .Z(n521) );
  and2 U532 ( .A1(w1), .A2(n469), .Z(n526) );
  and2 U533 ( .A1(a3), .A2(n470), .Z(n525) );
  or2 U534 ( .A1(n527), .A2(n528), .Z(n510) );
  and2 U535 ( .A1(n191), .A2(n196), .Z(n528) );
  inv1 U536 ( .I(n192), .ZN(n191) );
  and2 U537 ( .A1(n195), .A2(n192), .Z(n527) );
  or2 U538 ( .A1(n529), .A2(n530), .Z(n192) );
  or2 U539 ( .A1(n531), .A2(n532), .Z(n530) );
  and2 U540 ( .A1(n2), .A2(n465), .Z(n532) );
  and2 U541 ( .A1(x2), .A2(n466), .Z(n531) );
  or2 U542 ( .A1(n533), .A2(n534), .Z(n529) );
  and2 U543 ( .A1(d2), .A2(n469), .Z(n534) );
  and2 U544 ( .A1(h3), .A2(n470), .Z(n533) );
  inv1 U545 ( .I(n196), .ZN(n195) );
  or2 U546 ( .A1(n535), .A2(n536), .Z(n196) );
  or2 U547 ( .A1(n537), .A2(n538), .Z(n536) );
  and2 U548 ( .A1(o2), .A2(n465), .Z(n538) );
  and2 U550 ( .A1(y2), .A2(n466), .Z(n537) );
  or2 U552 ( .A1(n540), .A2(n541), .Z(n535) );
  and2 U553 ( .A1(e2), .A2(n469), .Z(n541) );
  and2 U555 ( .A1(i3), .A2(n470), .Z(n540) );
  inv1 U559 ( .I(i12), .ZN(b12) );
  or2 U560 ( .A1(n543), .A2(n544), .Z(i12) );
  or2 U561 ( .A1(n545), .A2(n546), .Z(n544) );
  and2 U562 ( .A1(u0), .A2(n446), .Z(n546) );
  and2 U563 ( .A1(k0), .A2(n447), .Z(n545) );
  or2 U564 ( .A1(n547), .A2(n548), .Z(n543) );
  and2 U565 ( .A1(f1), .A2(n450), .Z(n548) );
  and2 U566 ( .A1(q1), .A2(n451), .Z(n547) );
  or2 U567 ( .A1(n549), .A2(n550), .Z(a301) );
  and2 U568 ( .A1(n551), .A2(n216), .Z(n550) );
  inv1 U569 ( .I(q6), .ZN(n216) );
  and2 U570 ( .A1(n552), .A2(q6), .Z(n549) );
  and2 U571 ( .A1(n553), .A2(n554), .Z(n552) );
  or2 U572 ( .A1(n555), .A2(n426), .Z(n554) );
  inv1 U573 ( .I(n556), .ZN(n553) );
  and2 U574 ( .A1(n426), .A2(n555), .Z(n556) );
  or2 U575 ( .A1(n557), .A2(n558), .Z(n555) );
  and2 U576 ( .A1(n427), .A2(n207), .Z(n558) );
  inv1 U577 ( .I(n559), .ZN(n557) );
  or2 U578 ( .A1(n207), .A2(n427), .Z(n559) );
  or2 U579 ( .A1(n560), .A2(n561), .Z(n427) );
  inv1 U580 ( .I(n562), .ZN(n561) );
  or2 U581 ( .A1(n563), .A2(n564), .Z(n562) );
  and2 U582 ( .A1(n564), .A2(n563), .Z(n560) );
  inv1 U583 ( .I(n565), .ZN(n563) );
  or2 U584 ( .A1(n566), .A2(n567), .Z(n565) );
  and2 U585 ( .A1(n568), .A2(n131), .Z(n567) );
  and2 U586 ( .A1(n130), .A2(n551), .Z(n566) );
  or2 U587 ( .A1(n569), .A2(n570), .Z(n564) );
  and2 U588 ( .A1(n121), .A2(g12), .Z(n570) );
  and2 U589 ( .A1(n122), .A2(n127), .Z(n569) );
  inv1 U590 ( .I(g12), .ZN(n127) );
  or2 U591 ( .A1(n571), .A2(n572), .Z(g12) );
  or2 U592 ( .A1(n573), .A2(n574), .Z(n572) );
  and2 U593 ( .A1(w0), .A2(n446), .Z(n574) );
  and2 U594 ( .A1(m0), .A2(n447), .Z(n573) );
  or2 U595 ( .A1(n575), .A2(n576), .Z(n571) );
  and2 U596 ( .A1(h1), .A2(n450), .Z(n576) );
  and2 U597 ( .A1(s1), .A2(n451), .Z(n575) );
  and2 U598 ( .A1(n577), .A2(n578), .Z(n426) );
  or2 U599 ( .A1(n579), .A2(n580), .Z(n578) );
  inv1 U600 ( .I(n581), .ZN(n577) );
  and2 U601 ( .A1(n580), .A2(n579), .Z(n581) );
  inv1 U602 ( .I(n582), .ZN(n579) );
  or2 U603 ( .A1(n583), .A2(n584), .Z(n582) );
  and2 U604 ( .A1(k12), .A2(a12), .Z(n584) );
  and2 U605 ( .A1(j12), .A2(n146), .Z(n583) );
  inv1 U606 ( .I(k12), .ZN(n146) );
  or2 U607 ( .A1(n585), .A2(n586), .Z(k12) );
  or2 U608 ( .A1(n587), .A2(n588), .Z(n586) );
  and2 U609 ( .A1(o1), .A2(n589), .Z(n588) );
  and2 U610 ( .A1(d1), .A2(n6), .Z(n587) );
  or2 U611 ( .A1(n446), .A2(n590), .Z(n585) );
  and2 U612 ( .A1(i0), .A2(n447), .Z(n590) );
  or2 U613 ( .A1(n591), .A2(n592), .Z(n580) );
  and2 U614 ( .A1(m12), .A2(n151), .Z(n592) );
  inv1 U615 ( .I(l12), .ZN(n151) );
  and2 U616 ( .A1(l12), .A2(n154), .Z(n591) );
  inv1 U617 ( .I(m12), .ZN(n154) );
  or2 U618 ( .A1(n593), .A2(n594), .Z(m12) );
  or2 U619 ( .A1(n595), .A2(n596), .Z(n594) );
  and2 U620 ( .A1(r0), .A2(n446), .Z(n596) );
  and2 U621 ( .A1(g0), .A2(n447), .Z(n595) );
  or2 U622 ( .A1(n597), .A2(n598), .Z(n593) );
  and2 U623 ( .A1(b1), .A2(n450), .Z(n598) );
  and2 U624 ( .A1(m1), .A2(n451), .Z(n597) );
  or2 U625 ( .A1(n599), .A2(n600), .Z(l12) );
  or2 U626 ( .A1(n601), .A2(n602), .Z(n600) );
  and2 U627 ( .A1(s0), .A2(n446), .Z(n602) );
  and2 U628 ( .A1(h0), .A2(n447), .Z(n601) );
  or2 U629 ( .A1(n603), .A2(n604), .Z(n599) );
  and2 U630 ( .A1(c1), .A2(n450), .Z(n604) );
  and2 U631 ( .A1(n1), .A2(n451), .Z(n603) );
  and2 U632 ( .A1(n605), .A2(n606), .Z(a13) );
  or2 U633 ( .A1(n607), .A2(n551), .Z(n606) );
  inv1 U634 ( .I(n608), .ZN(n607) );
  or2 U635 ( .A1(n568), .A2(n608), .Z(n605) );
  or2 U636 ( .A1(p6), .A2(n609), .Z(n608) );
  and2 U637 ( .A1(n610), .A2(n611), .Z(n609) );
  or2 U638 ( .A1(n612), .A2(n207), .Z(n611) );
  inv1 U639 ( .I(n613), .ZN(n610) );
  and2 U640 ( .A1(n207), .A2(n612), .Z(n613) );
  or2 U641 ( .A1(n614), .A2(n615), .Z(n612) );
  and2 U642 ( .A1(n130), .A2(n122), .Z(n615) );
  inv1 U643 ( .I(n131), .ZN(n130) );
  and2 U644 ( .A1(n121), .A2(n131), .Z(n614) );
  or2 U645 ( .A1(n616), .A2(n617), .Z(n131) );
  or2 U646 ( .A1(n618), .A2(n619), .Z(n617) );
  and2 U647 ( .A1(p0), .A2(n446), .Z(n619) );
  and2 U648 ( .A1(e0), .A2(n447), .Z(n618) );
  or2 U649 ( .A1(n620), .A2(n621), .Z(n616) );
  and2 U650 ( .A1(z0), .A2(n450), .Z(n621) );
  and2 U651 ( .A1(k1), .A2(n451), .Z(n620) );
  inv1 U652 ( .I(n122), .ZN(n121) );
  or2 U653 ( .A1(l6), .A2(n122), .Z(n207) );
  or2 U654 ( .A1(n622), .A2(n623), .Z(n122) );
  or2 U655 ( .A1(n624), .A2(n625), .Z(n623) );
  and2 U656 ( .A1(x0), .A2(n446), .Z(n625) );
  and2 U657 ( .A1(n0), .A2(n447), .Z(n624) );
  or2 U658 ( .A1(n626), .A2(n627), .Z(n622) );
  and2 U659 ( .A1(i1), .A2(n450), .Z(n627) );
  and2 U660 ( .A1(t1), .A2(n451), .Z(n626) );
  inv1 U661 ( .I(n551), .ZN(n568) );
  or2 U662 ( .A1(n628), .A2(n629), .Z(n551) );
  or2 U663 ( .A1(n630), .A2(n631), .Z(n629) );
  and2 U664 ( .A1(y0), .A2(n446), .Z(n631) );
  and2 U665 ( .A1(o0), .A2(n447), .Z(n630) );
  or2 U666 ( .A1(n632), .A2(n633), .Z(n628) );
  and2 U667 ( .A1(j1), .A2(n450), .Z(n633) );
  and2 U668 ( .A1(u1), .A2(n451), .Z(n632) );
  inv1 U669 ( .I(j12), .ZN(a12) );
  or2 U670 ( .A1(n634), .A2(n635), .Z(j12) );
  or2 U671 ( .A1(n636), .A2(n637), .Z(n635) );
  and2 U672 ( .A1(t0), .A2(n446), .Z(n637) );
  and2 U673 ( .A1(n589), .A2(n6), .Z(n446) );
  and2 U674 ( .A1(j0), .A2(n447), .Z(n636) );
  and2 U675 ( .A1(n638), .A2(k6), .Z(n447) );
  or2 U676 ( .A1(n639), .A2(n640), .Z(n634) );
  and2 U677 ( .A1(e1), .A2(n450), .Z(n640) );
  and2 U678 ( .A1(k6), .A2(n6), .Z(n450) );
  and2 U679 ( .A1(p1), .A2(n451), .Z(n639) );
  and2 U680 ( .A1(n638), .A2(n589), .Z(n451) );
  inv1 U681 ( .I(k6), .ZN(n589) );
  inv1 U682 ( .I(n6), .ZN(n638) );
  and2 U683 ( .A1(n379), .A2(n34), .Z(n391) );
  and2 U684 ( .A1(n378), .A2(n87), .Z(n392) );
  or2 U685 ( .A1(n499), .A2(n500), .Z(n495) );
  or2 U686 ( .A1(n359), .A2(n360), .Z(n358) );
  and2f U687 ( .A1(n363), .A2(n364), .Z(n359) );
  and2f U688 ( .A1(n351), .A2(n352), .Z(n347) );
  or2f U689 ( .A1(n353), .A2(n354), .Z(n352) );
  or2f U690 ( .A1(n463), .A2(n464), .Z(n462) );
  or2f U691 ( .A1(n467), .A2(n468), .Z(n461) );
  and2f U692 ( .A1(n410), .A2(n174), .Z(n408) );
  or2f U693 ( .A1(n495), .A2(n496), .Z(n174) );
  inv1f U694 ( .I(n171), .ZN(x11) );
  or2f U695 ( .A1(n461), .A2(n462), .Z(n171) );
  and2f U696 ( .A1(n379), .A2(n38), .Z(n393) );
  inv1f U697 ( .I(n379), .ZN(n378) );
  inv1f U698 ( .I(n7), .ZN(n542) );
  and2f U699 ( .A1(u2), .A2(n466), .Z(n463) );
  and2f U700 ( .A1(v2), .A2(n466), .Z(n497) );
  and2f U701 ( .A1(n408), .A2(n409), .Z(n379) );
  and2f U702 ( .A1(x11), .A2(d0), .Z(n409) );
  and2f U703 ( .A1(k2), .A2(n465), .Z(n464) );
  and2f U704 ( .A1(l2), .A2(n465), .Z(n498) );
  and2f U705 ( .A1(m7), .A2(n7), .Z(n465) );
  and2f U706 ( .A1(e3), .A2(n470), .Z(n467) );
  and2f U707 ( .A1(f3), .A2(n470), .Z(n499) );
  and2f U708 ( .A1(n542), .A2(n539), .Z(n470) );
  and2f U709 ( .A1(n539), .A2(n7), .Z(n466) );
  inv1f U710 ( .I(m7), .ZN(n539) );
  and2f U711 ( .A1(a2), .A2(n469), .Z(n468) );
  and2f U712 ( .A1(b2), .A2(n469), .Z(n500) );
  and2f U713 ( .A1(n542), .A2(m7), .Z(n469) );
  or2 U714 ( .A1(n380), .A2(n381), .Z(n373) );
  and2 U715 ( .A1(n383), .A2(n384), .Z(n380) );
  and2 U716 ( .A1(n375), .A2(c12), .Z(n371) );
  or2 U717 ( .A1(n373), .A2(n374), .Z(n375) );
  or2 U718 ( .A1(n365), .A2(n366), .Z(n364) );
  or2 U719 ( .A1(n334), .A2(n335), .Z(n333) );
  or2 U720 ( .A1(n322), .A2(n323), .Z(f13) );
  and2 U721 ( .A1(n326), .A2(n327), .Z(n322) );
  and2f U722 ( .A1(n345), .A2(n346), .Z(n342) );
  or2f U723 ( .A1(n347), .A2(n348), .Z(n346) );
  and2f U724 ( .A1(n342), .A2(n340), .Z(n336) );
  and2f U725 ( .A1(n369), .A2(n370), .Z(n365) );
  or2f U726 ( .A1(n371), .A2(n372), .Z(n370) );
  and2f U727 ( .A1(n357), .A2(n358), .Z(n353) );
  or2f U728 ( .A1(n328), .A2(n329), .Z(n327) );
  or2f U729 ( .A1(n393), .A2(n394), .Z(n387) );
  and2f U730 ( .A1(n378), .A2(n73), .Z(n394) );
  and2f U731 ( .A1(n332), .A2(n333), .Z(n328) );
endmodule

