
module count ( j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, s, r, 
        q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, z0, y0, x0, w0, v0, 
        u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0 );
  input j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, s, r, q, p,
         o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0;
  wire   n67, n68, n69, n74, n75, n76, n77, n83, n84, n85, n86, n87, n88, n89,
         n90, n93, n94, n95, n96, n97, n103, n104, n105, n106, n107, n108,
         n109, n110, n113, n114, n115, n116, n117, n121, n122, n123, n124,
         n128, n129, n130, n131, n138, n139, n140, n141, n142, n143, n144,
         n145, n148, n149, n150, n151, n152, n155, n158, n159, n160, n161,
         n162, n163, n164, n165, n168, n169, n170, n171, n172, n176, n177,
         n178, n179, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n259, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271;

  or2f U34 ( .A1(s), .A2(n69), .Z(n68) );
  or2f U43 ( .A1(s), .A2(n77), .Z(n76) );
  or2f U53 ( .A1(n84), .A2(n85), .Z(u0) );
  or2f U54 ( .A1(s), .A2(n86), .Z(n85) );
  and2f U55 ( .A1(n87), .A2(q), .Z(n86) );
  and2f U56 ( .A1(n88), .A2(n89), .Z(n87) );
  or2f U64 ( .A1(s), .A2(n96), .Z(n95) );
  and2f U65 ( .A1(q), .A2(n97), .Z(n96) );
  or2f U75 ( .A1(n104), .A2(n105), .Z(s0) );
  or2f U76 ( .A1(n106), .A2(s), .Z(n105) );
  and2f U77 ( .A1(n107), .A2(q), .Z(n106) );
  and2f U78 ( .A1(n108), .A2(n109), .Z(n107) );
  or2f U86 ( .A1(s), .A2(n116), .Z(n115) );
  and2f U87 ( .A1(q), .A2(n117), .Z(n116) );
  and2 U167 ( .A1(h0), .A2(n235), .Z(n236) );
  and2 U168 ( .A1(n254), .A2(q), .Z(n246) );
  inv1 U170 ( .I(n197), .ZN(n187) );
  inv1 U171 ( .I(n230), .ZN(n227) );
  and2 U172 ( .A1(q), .A2(n243), .Z(n238) );
  inv1 U173 ( .I(n223), .ZN(n202) );
  and2 U174 ( .A1(i0), .A2(n243), .Z(n244) );
  and2 U175 ( .A1(a0), .A2(n223), .Z(n206) );
  and2 U176 ( .A1(v), .A2(n197), .Z(n189) );
  or2 U178 ( .A1(n197), .A2(v), .Z(n193) );
  or2 U179 ( .A1(n197), .A2(v), .Z(n191) );
  or2f U183 ( .A1(u), .A2(r), .Z(n197) );
  or2f U191 ( .A1(v), .A2(w), .Z(n198) );
  or2f U197 ( .A1(n198), .A2(n197), .Z(n200) );
  or2f U201 ( .A1(n261), .A2(n200), .Z(n223) );
  or2f U210 ( .A1(n209), .A2(n208), .Z(n117) );
  and2f U211 ( .A1(n110), .A2(n210), .Z(n211) );
  or2f U217 ( .A1(n219), .A2(d0), .Z(n216) );
  or2f U220 ( .A1(n215), .A2(n214), .Z(n97) );
  and2f U221 ( .A1(n216), .A2(n90), .Z(n217) );
  and2f U227 ( .A1(f0), .A2(n220), .Z(n228) );
  or2f U228 ( .A1(n222), .A2(n221), .Z(n224) );
  or2f U229 ( .A1(n224), .A2(n223), .Z(n226) );
  or2f U232 ( .A1(n228), .A2(n227), .Z(n229) );
  and2f U233 ( .A1(q), .A2(n229), .Z(n77) );
  or2f U234 ( .A1(n185), .A2(n226), .Z(n235) );
  inv1f U235 ( .I(n231), .ZN(n232) );
  and2f U236 ( .A1(n235), .A2(n232), .Z(n233) );
  or2f U237 ( .A1(n233), .A2(n186), .Z(n234) );
  inv1f U238 ( .I(n234), .ZN(n69) );
  or2f U239 ( .A1(n270), .A2(n226), .Z(n243) );
  inv1f U240 ( .I(n236), .ZN(n237) );
  and2f U241 ( .A1(n238), .A2(n237), .Z(n240) );
  or2f U243 ( .A1(n240), .A2(n239), .Z(n241) );
  inv1f U244 ( .I(n241), .ZN(n242) );
  inv1f U247 ( .I(n244), .ZN(n245) );
  and2f U248 ( .A1(n246), .A2(n245), .Z(n248) );
  or2f U250 ( .A1(n248), .A2(n247), .Z(n249) );
  inv1f U251 ( .I(n249), .ZN(n250) );
  and2f U256 ( .A1(n254), .A2(n253), .Z(n252) );
  and2f U258 ( .A1(n256), .A2(n255), .Z(n257) );
  or2 U164 ( .A1(d0), .A2(e0), .Z(n222) );
  or2f U165 ( .A1(n219), .A2(n222), .Z(n220) );
  or2 U166 ( .A1(n254), .A2(n253), .Z(n255) );
  or2f U169 ( .A1(n226), .A2(n271), .Z(n254) );
  inv1 U177 ( .I(n252), .ZN(n256) );
  or2f U180 ( .A1(n265), .A2(n223), .Z(n230) );
  or2 U181 ( .A1(n200), .A2(n199), .Z(n201) );
  inv1 U182 ( .I(n267), .ZN(n266) );
  inv1 U184 ( .I(a0), .ZN(n268) );
  inv1 U185 ( .I(n221), .ZN(n269) );
  and2 U186 ( .A1(g0), .A2(n230), .Z(n231) );
  or2 U187 ( .A1(n183), .A2(n194), .Z(n152) );
  and2 U188 ( .A1(n142), .A2(q), .Z(n141) );
  and2 U189 ( .A1(n143), .A2(n144), .Z(n142) );
  or2 U190 ( .A1(n196), .A2(n145), .Z(n144) );
  or2 U192 ( .A1(n183), .A2(y), .Z(n143) );
  or2 U193 ( .A1(n203), .A2(n202), .Z(n204) );
  or2 U194 ( .A1(n210), .A2(n110), .Z(n109) );
  inv1 U195 ( .I(n211), .ZN(n108) );
  or2 U196 ( .A1(n216), .A2(n90), .Z(n89) );
  inv1 U198 ( .I(n217), .ZN(n88) );
  or2 U199 ( .A1(n114), .A2(n115), .Z(r0) );
  or2 U200 ( .A1(n94), .A2(n95), .Z(t0) );
  or2 U202 ( .A1(n75), .A2(n76), .Z(v0) );
  or2 U203 ( .A1(n67), .A2(n68), .Z(w0) );
  or2 U204 ( .A1(n242), .A2(s), .Z(x0) );
  and2 U205 ( .A1(c), .A2(n186), .Z(n239) );
  or2 U206 ( .A1(n250), .A2(s), .Z(y0) );
  and2 U207 ( .A1(b), .A2(n186), .Z(n247) );
  and2 U208 ( .A1(n262), .A2(n263), .Z(z0) );
  inv1 U209 ( .I(n213), .ZN(n205) );
  or2f U212 ( .A1(n198), .A2(n197), .Z(n195) );
  or2f U213 ( .A1(z), .A2(n199), .Z(n261) );
  or2 U214 ( .A1(x), .A2(y), .Z(n199) );
  or2 U215 ( .A1(n257), .A2(n264), .Z(n262) );
  or2 U216 ( .A1(s), .A2(n259), .Z(n263) );
  or2 U218 ( .A1(n186), .A2(s), .Z(n264) );
  or2 U219 ( .A1(n219), .A2(d0), .Z(n218) );
  or2 U222 ( .A1(n213), .A2(b0), .Z(n212) );
  or2 U223 ( .A1(n224), .A2(n225), .Z(n265) );
  or2f U224 ( .A1(n213), .A2(b0), .Z(n210) );
  inv1 U225 ( .I(n212), .ZN(n209) );
  or2f U226 ( .A1(n223), .A2(n266), .Z(n219) );
  inv1 U230 ( .I(n218), .ZN(n215) );
  and2f U231 ( .A1(n268), .A2(n269), .Z(n267) );
  or2 U242 ( .A1(b0), .A2(c0), .Z(n221) );
  and2 U245 ( .A1(b0), .A2(n213), .Z(n208) );
  or2f U246 ( .A1(n223), .A2(a0), .Z(n213) );
  and2 U249 ( .A1(d0), .A2(n219), .Z(n214) );
  or2f U252 ( .A1(n185), .A2(h0), .Z(n270) );
  or2f U253 ( .A1(n270), .A2(i0), .Z(n271) );
  or2 U254 ( .A1(a0), .A2(f0), .Z(n225) );
  and2 U255 ( .A1(q), .A2(n188), .Z(n179) );
  or2 U257 ( .A1(n187), .A2(n181), .Z(n188) );
  and2 U259 ( .A1(u), .A2(r), .Z(n181) );
  or2 U260 ( .A1(q), .A2(p), .Z(n182) );
  and2 U261 ( .A1(q), .A2(n172), .Z(n171) );
  or2 U262 ( .A1(n190), .A2(n189), .Z(n172) );
  inv1 U263 ( .I(n191), .ZN(n190) );
  or2 U264 ( .A1(q), .A2(o), .Z(n176) );
  and2 U265 ( .A1(n162), .A2(q), .Z(n161) );
  and2 U266 ( .A1(n163), .A2(n164), .Z(n162) );
  or2 U267 ( .A1(n193), .A2(n165), .Z(n164) );
  inv1 U268 ( .I(n192), .ZN(n163) );
  or2 U269 ( .A1(q), .A2(n), .Z(n168) );
  and2 U270 ( .A1(q), .A2(n152), .Z(n151) );
  and2 U271 ( .A1(x), .A2(n195), .Z(n194) );
  or2 U272 ( .A1(q), .A2(m), .Z(n158) );
  or2 U273 ( .A1(q), .A2(l), .Z(n148) );
  and2 U274 ( .A1(q), .A2(n204), .Z(n131) );
  and2 U275 ( .A1(z), .A2(n201), .Z(n203) );
  or2 U276 ( .A1(q), .A2(k), .Z(n138) );
  inv1 U277 ( .I(q), .ZN(n186) );
  inv1 U278 ( .I(a), .ZN(n251) );
  and2 U279 ( .A1(n165), .A2(n191), .Z(n192) );
  inv1 U280 ( .I(w), .ZN(n165) );
  or2 U281 ( .A1(n195), .A2(x), .Z(n196) );
  inv1 U282 ( .I(y), .ZN(n145) );
  and2 U283 ( .A1(n184), .A2(n155), .Z(n183) );
  inv1 U284 ( .I(x), .ZN(n155) );
  inv1 U285 ( .I(n195), .ZN(n184) );
  inv1 U286 ( .I(c0), .ZN(n110) );
  inv1 U287 ( .I(e0), .ZN(n90) );
  or2 U288 ( .A1(g0), .A2(n225), .Z(n185) );
  inv1 U289 ( .I(j0), .ZN(n253) );
  and2 U290 ( .A1(n207), .A2(q), .Z(n124) );
  or2 U291 ( .A1(n206), .A2(n205), .Z(n207) );
  inv1 U292 ( .I(n182), .ZN(n177) );
  or2 U293 ( .A1(s), .A2(n179), .Z(n178) );
  inv1 U294 ( .I(n176), .ZN(n169) );
  or2 U295 ( .A1(s), .A2(n171), .Z(n170) );
  inv1 U296 ( .I(n168), .ZN(n159) );
  or2 U297 ( .A1(s), .A2(n161), .Z(n160) );
  inv1 U298 ( .I(n158), .ZN(n149) );
  or2 U299 ( .A1(s), .A2(n151), .Z(n150) );
  inv1 U300 ( .I(n148), .ZN(n139) );
  or2 U301 ( .A1(s), .A2(n141), .Z(n140) );
  inv1 U302 ( .I(n138), .ZN(n129) );
  or2 U303 ( .A1(s), .A2(n131), .Z(n130) );
  or2 U304 ( .A1(n122), .A2(n123), .Z(q0) );
  inv1 U305 ( .I(n128), .ZN(n122) );
  or2 U306 ( .A1(s), .A2(n124), .Z(n123) );
  or2 U307 ( .A1(q), .A2(j), .Z(n128) );
  inv1 U308 ( .I(n121), .ZN(n114) );
  or2 U309 ( .A1(q), .A2(i), .Z(n121) );
  inv1 U310 ( .I(n113), .ZN(n104) );
  or2 U311 ( .A1(q), .A2(h), .Z(n113) );
  inv1 U312 ( .I(n103), .ZN(n94) );
  or2 U313 ( .A1(q), .A2(g), .Z(n103) );
  inv1 U314 ( .I(n93), .ZN(n84) );
  or2 U315 ( .A1(q), .A2(f), .Z(n93) );
  inv1 U316 ( .I(n83), .ZN(n75) );
  or2 U317 ( .A1(q), .A2(e), .Z(n83) );
  inv1 U318 ( .I(n74), .ZN(n67) );
  or2 U319 ( .A1(q), .A2(d), .Z(n74) );
  or2 U320 ( .A1(q), .A2(n251), .Z(n259) );
  or2 U321 ( .A1(n177), .A2(n178), .Z(k0) );
  or2 U322 ( .A1(n169), .A2(n170), .Z(l0) );
  or2 U323 ( .A1(n159), .A2(n160), .Z(m0) );
  or2 U324 ( .A1(n149), .A2(n150), .Z(n0) );
  or2 U325 ( .A1(n139), .A2(n140), .Z(o0) );
  or2 U326 ( .A1(n129), .A2(n130), .Z(p0) );
endmodule

