
module x4 ( v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, g2, f2, 
        e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, 
        m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, 
        u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, i0, h0, g0, f0, e0, d0, c0, 
        b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, i, h, g, b, a, 
        o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4, x4, 
        w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4, h4, g4, f4, 
        e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, o3, n3, 
        m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, y2, x2, w2 );
  input v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, g2, f2, e2,
         d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1,
         m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, w0,
         v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, i0, h0, g0, f0, e0,
         d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, i, h,
         g, b, a;
  output o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4, y4,
         x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4, h4,
         g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3,
         p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2,
         y2, x2, w2;
  wire   n13, n14, n15, n16, n18, n23, n24, n25, n35, n73, n74, n77, n78, n92,
         n93, n94, n95, n96, n97, n102, n103, n104, n105, n106, n165, n166,
         n167, n169, n170, n171, n172, n173, n178, n179, n180, n209, n210,
         n211, n212, n213, n214, n216, n217, n222, n223, n224, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n244, n250, n251, n252, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n279, n280, n281,
         n284, n285, n286, n287, n288, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n520, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544;

  and2 U6 ( .A1(n13), .A2(n14), .Z(z3) );
  or2 U7 ( .A1(p0), .A2(n541), .Z(n14) );
  and2 U8 ( .A1(n16), .A2(n307), .Z(n13) );
  or2 U9 ( .A1(n540), .A2(g1), .Z(n16) );
  inv1 U10 ( .I(i1), .ZN(z2) );
  and2 U16 ( .A1(n23), .A2(n24), .Z(y3) );
  or2 U17 ( .A1(o0), .A2(n541), .Z(n24) );
  and2 U18 ( .A1(n25), .A2(n307), .Z(n23) );
  or2 U19 ( .A1(n18), .A2(f1), .Z(n25) );
  inv1 U20 ( .I(h1), .ZN(y2) );
  inv1 U27 ( .I(g1), .ZN(x2) );
  and2 U37 ( .A1(i0), .A2(v2), .Z(n35) );
  inv1 U38 ( .I(f1), .ZN(w2) );
  and2 U51 ( .A1(a1), .A2(n524), .Z(u3) );
  and2 U57 ( .A1(z0), .A2(n524), .Z(t3) );
  and2 U63 ( .A1(y0), .A2(n524), .Z(s3) );
  and2 U69 ( .A1(x0), .A2(n524), .Z(r3) );
  and2 U75 ( .A1(w0), .A2(n524), .Z(q3) );
  and2 U81 ( .A1(v0), .A2(n524), .Z(p3) );
  and2 U82 ( .A1(n73), .A2(n524), .Z(o5) );
  and2 U85 ( .A1(n77), .A2(v2), .Z(n74) );
  inv1 U86 ( .I(n78), .ZN(n77) );
  or2 U87 ( .A1(f0), .A2(g0), .Z(n78) );
  and2 U93 ( .A1(a), .A2(n524), .Z(o3) );
  and2 U102 ( .A1(b), .A2(n524), .Z(n3) );
  and2 U103 ( .A1(n92), .A2(n307), .Z(m5) );
  or2 U104 ( .A1(n93), .A2(n94), .Z(n92) );
  and2 U105 ( .A1(n95), .A2(n96), .Z(n94) );
  and2 U106 ( .A1(t2), .A2(n97), .Z(n93) );
  inv1 U107 ( .I(n95), .ZN(n97) );
  and2 U108 ( .A1(l1), .A2(s2), .Z(n95) );
  and2 U114 ( .A1(t0), .A2(n102), .Z(m3) );
  and2 U115 ( .A1(n103), .A2(n524), .Z(l5) );
  or2 U116 ( .A1(n104), .A2(n105), .Z(n103) );
  and2 U117 ( .A1(b1), .A2(n106), .Z(n105) );
  and2 U118 ( .A1(n1), .A2(n305), .Z(n104) );
  and2 U124 ( .A1(s0), .A2(n102), .Z(l3) );
  and2 U136 ( .A1(r0), .A2(n102), .Z(k3) );
  and2 U150 ( .A1(q0), .A2(n102), .Z(j3) );
  and2 U165 ( .A1(p0), .A2(n102), .Z(i3) );
  and2 U179 ( .A1(o0), .A2(n102), .Z(h3) );
  or2 U187 ( .A1(n165), .A2(n166), .Z(g4) );
  and2 U188 ( .A1(n167), .A2(i), .Z(n166) );
  and2 U189 ( .A1(n518), .A2(g0), .Z(n167) );
  or2 U191 ( .A1(n171), .A2(n172), .Z(n170) );
  and2 U192 ( .A1(n1), .A2(n106), .Z(n172) );
  and2 U193 ( .A1(n534), .A2(n173), .Z(n171) );
  inv1 U194 ( .I(o1), .ZN(n173) );
  or2 U199 ( .A1(n178), .A2(n179), .Z(g3) );
  and2 U200 ( .A1(n180), .A2(n524), .Z(n179) );
  and2 U201 ( .A1(n0), .A2(n102), .Z(n178) );
  and2 U202 ( .A1(n524), .A2(n307), .Z(n102) );
  or2 U233 ( .A1(n209), .A2(n180), .Z(e4) );
  and2 U234 ( .A1(l1), .A2(n307), .Z(n209) );
  or2 U235 ( .A1(n210), .A2(n180), .Z(e3) );
  inv1 U236 ( .I(n211), .ZN(n180) );
  or2 U237 ( .A1(n212), .A2(n213), .Z(n211) );
  or2 U238 ( .A1(n522), .A2(n214), .Z(n213) );
  or2 U239 ( .A1(n523), .A2(c1), .Z(n214) );
  or2 U240 ( .A1(n216), .A2(n217), .Z(n212) );
  and2 U241 ( .A1(l0), .A2(n307), .Z(n210) );
  and2 U251 ( .A1(n222), .A2(n223), .Z(d4) );
  or2 U252 ( .A1(t0), .A2(n541), .Z(n223) );
  and2 U253 ( .A1(n224), .A2(n307), .Z(n222) );
  or2 U254 ( .A1(n18), .A2(k1), .Z(n224) );
  and2 U263 ( .A1(n230), .A2(n231), .Z(c4) );
  or2 U264 ( .A1(s0), .A2(n541), .Z(n231) );
  and2 U265 ( .A1(n232), .A2(n307), .Z(n230) );
  or2 U266 ( .A1(n18), .A2(j1), .Z(n232) );
  and2 U267 ( .A1(n233), .A2(n524), .Z(c3) );
  or2 U268 ( .A1(n234), .A2(n235), .Z(n233) );
  and2 U269 ( .A1(s2), .A2(n236), .Z(n235) );
  and2 U270 ( .A1(n237), .A2(n538), .Z(n234) );
  or2 U273 ( .A1(n520), .A2(n240), .Z(n239) );
  or2 U278 ( .A1(p2), .A2(o2), .Z(n217) );
  inv1 U279 ( .I(n242), .ZN(n241) );
  or2 U280 ( .A1(i), .A2(q2), .Z(n242) );
  or2 U282 ( .A1(h0), .A2(n96), .Z(n244) );
  inv1 U283 ( .I(t2), .ZN(n96) );
  and2 U290 ( .A1(n250), .A2(n251), .Z(b4) );
  or2 U291 ( .A1(r0), .A2(n541), .Z(n251) );
  and2 U292 ( .A1(n252), .A2(n307), .Z(n250) );
  or2 U293 ( .A1(n539), .A2(i1), .Z(n252) );
  inv1 U294 ( .I(k1), .ZN(b3) );
  and2 U320 ( .A1(n262), .A2(n263), .Z(a4) );
  or2 U321 ( .A1(q0), .A2(n541), .Z(n263) );
  and2 U322 ( .A1(n264), .A2(n307), .Z(n262) );
  or2 U324 ( .A1(n540), .A2(h1), .Z(n264) );
  or2 U332 ( .A1(r2), .A2(q2), .Z(n216) );
  inv1 U333 ( .I(j1), .ZN(a3) );
  or2 U334 ( .A1(n273), .A2(n269), .Z(n268) );
  inv1 U335 ( .I(n268), .ZN(n274) );
  inv1 U336 ( .I(m2), .ZN(n269) );
  or2 U342 ( .A1(h), .A2(i), .Z(n276) );
  inv1 U347 ( .I(u0), .ZN(n281) );
  buf0 U348 ( .I(n517), .Z(x3) );
  or2 U352 ( .A1(n531), .A2(g), .Z(n287) );
  or2 U356 ( .A1(n351), .A2(n352), .Z(n290) );
  or2 U360 ( .A1(n293), .A2(n294), .Z(n299) );
  or2 U364 ( .A1(n314), .A2(n325), .Z(n296) );
  inv1 U370 ( .I(n303), .ZN(n334) );
  and2 U372 ( .A1(e1), .A2(n306), .Z(n305) );
  inv1 U373 ( .I(n534), .ZN(n106) );
  inv1 U375 ( .I(c1), .ZN(n307) );
  inv1 U379 ( .I(e1), .ZN(n523) );
  inv1 U381 ( .I(r2), .ZN(n520) );
  or2 U383 ( .A1(n530), .A2(t2), .Z(n310) );
  and2 U384 ( .A1(n244), .A2(n310), .Z(n237) );
  inv1 U387 ( .I(i0), .ZN(n524) );
  inv1 U388 ( .I(h), .ZN(n346) );
  or2 U389 ( .A1(n350), .A2(g), .Z(n327) );
  inv1 U390 ( .I(n287), .ZN(n311) );
  and2 U391 ( .A1(n346), .A2(n311), .Z(n312) );
  or2 U396 ( .A1(n342), .A2(n527), .Z(n328) );
  or2 U397 ( .A1(n312), .A2(n328), .Z(n313) );
  and2 U398 ( .A1(n524), .A2(n313), .Z(n169) );
  or2 U400 ( .A1(n315), .A2(i0), .Z(n363) );
  inv1 U401 ( .I(n363), .ZN(n518) );
  and2 U402 ( .A1(n538), .A2(n342), .Z(n316) );
  or2 U403 ( .A1(n316), .A2(n74), .Z(n73) );
  and2 U405 ( .A1(g), .A2(m1), .Z(n318) );
  or2 U406 ( .A1(n319), .A2(n318), .Z(n320) );
  and2 U408 ( .A1(h), .A2(m1), .Z(n322) );
  and2 U409 ( .A1(i), .A2(m1), .Z(n321) );
  inv1 U411 ( .I(f0), .ZN(n325) );
  or2 U412 ( .A1(n334), .A2(k0), .Z(n326) );
  and2 U413 ( .A1(n307), .A2(n326), .Z(d3) );
  or2 U414 ( .A1(h), .A2(i), .Z(n352) );
  or2 U417 ( .A1(n432), .A2(n328), .Z(n331) );
  inv1 U418 ( .I(n342), .ZN(n329) );
  or2 U419 ( .A1(n329), .A2(m0), .Z(n330) );
  and2 U420 ( .A1(n331), .A2(n330), .Z(n332) );
  or2 U421 ( .A1(n332), .A2(i0), .Z(f3) );
  or2 U422 ( .A1(i0), .A2(n538), .Z(n333) );
  or2 U423 ( .A1(n334), .A2(n333), .Z(v3) );
  and2 U424 ( .A1(n362), .A2(n35), .Z(n338) );
  and2 U425 ( .A1(n527), .A2(n335), .Z(n337) );
  and2 U426 ( .A1(n338), .A2(n337), .Z(w3) );
  inv1 U429 ( .I(n272), .ZN(n343) );
  or2 U430 ( .A1(e1), .A2(d1), .Z(n340) );
  and2 U435 ( .A1(n524), .A2(n342), .Z(n349) );
  inv1 U436 ( .I(g), .ZN(n344) );
  and2 U437 ( .A1(n344), .A2(n343), .Z(n345) );
  and2 U438 ( .A1(n346), .A2(n345), .Z(n347) );
  and2 U440 ( .A1(n349), .A2(n348), .Z(f4) );
  or2 U442 ( .A1(n531), .A2(g), .Z(n351) );
  inv1 U447 ( .I(p1), .ZN(n356) );
  or2 U448 ( .A1(n106), .A2(n356), .Z(n358) );
  or2 U449 ( .A1(n305), .A2(o1), .Z(n357) );
  and2 U450 ( .A1(n358), .A2(n357), .Z(n359) );
  or2 U451 ( .A1(n359), .A2(i0), .Z(n360) );
  or2 U452 ( .A1(n532), .A2(n360), .Z(h4) );
  or2 U457 ( .A1(n294), .A2(n315), .Z(n433) );
  or2 U461 ( .A1(n366), .A2(n365), .Z(n370) );
  or2 U462 ( .A1(n106), .A2(i0), .Z(n367) );
  and2 U464 ( .A1(q1), .A2(n308), .Z(n369) );
  or2 U465 ( .A1(n370), .A2(n369), .Z(i4) );
  or2 U468 ( .A1(n372), .A2(n371), .Z(n374) );
  and2 U469 ( .A1(r1), .A2(n308), .Z(n373) );
  or2 U470 ( .A1(n374), .A2(n373), .Z(j4) );
  and2 U472 ( .A1(m), .A2(n387), .Z(n375) );
  and2 U474 ( .A1(s1), .A2(n526), .Z(n377) );
  or2 U475 ( .A1(n378), .A2(n377), .Z(k4) );
  and2 U477 ( .A1(n), .A2(n387), .Z(n379) );
  or2 U480 ( .A1(n382), .A2(n381), .Z(l4) );
  or2 U483 ( .A1(n384), .A2(n383), .Z(n386) );
  or2 U485 ( .A1(n386), .A2(n385), .Z(m4) );
  or2 U490 ( .A1(n391), .A2(n390), .Z(n4) );
  and2 U492 ( .A1(q), .A2(n387), .Z(n392) );
  and2 U494 ( .A1(w1), .A2(n543), .Z(n394) );
  or2 U495 ( .A1(n395), .A2(n394), .Z(o4) );
  or2 U498 ( .A1(n397), .A2(n396), .Z(n399) );
  and2 U499 ( .A1(x1), .A2(n526), .Z(n398) );
  or2 U500 ( .A1(n399), .A2(n398), .Z(p4) );
  and2 U501 ( .A1(x1), .A2(n544), .Z(n401) );
  or2 U505 ( .A1(n403), .A2(n402), .Z(q4) );
  and2 U506 ( .A1(n457), .A2(y1), .Z(n405) );
  and2 U507 ( .A1(t), .A2(n387), .Z(n404) );
  or2 U510 ( .A1(n407), .A2(n406), .Z(r4) );
  or2 U513 ( .A1(n410), .A2(n409), .Z(n412) );
  and2 U514 ( .A1(a2), .A2(n543), .Z(n411) );
  or2 U515 ( .A1(n412), .A2(n411), .Z(s4) );
  and2 U522 ( .A1(b2), .A2(n526), .Z(n418) );
  or2 U523 ( .A1(n419), .A2(n418), .Z(t4) );
  and2 U524 ( .A1(n408), .A2(b2), .Z(n421) );
  and2 U527 ( .A1(c2), .A2(n308), .Z(n422) );
  or2 U528 ( .A1(n423), .A2(n422), .Z(u4) );
  and2 U530 ( .A1(x), .A2(n456), .Z(n424) );
  and2 U532 ( .A1(d2), .A2(n308), .Z(n426) );
  or2 U533 ( .A1(n427), .A2(n426), .Z(v4) );
  and2 U534 ( .A1(n408), .A2(d2), .Z(n429) );
  and2 U537 ( .A1(e2), .A2(n543), .Z(n430) );
  or2 U538 ( .A1(n431), .A2(n430), .Z(w4) );
  or2 U543 ( .A1(n436), .A2(n435), .Z(n438) );
  or2 U545 ( .A1(n438), .A2(n437), .Z(x4) );
  or2 U550 ( .A1(n442), .A2(n441), .Z(y4) );
  or2 U555 ( .A1(n446), .A2(n445), .Z(z4) );
  or2 U560 ( .A1(n450), .A2(n449), .Z(a5) );
  and2 U562 ( .A1(d0), .A2(n451), .Z(n452) );
  or2 U565 ( .A1(n455), .A2(n454), .Z(b5) );
  and2 U566 ( .A1(e0), .A2(n456), .Z(n459) );
  and2 U567 ( .A1(j2), .A2(n301), .Z(n458) );
  or2 U568 ( .A1(n459), .A2(n458), .Z(c5) );
  inv1 U569 ( .I(k2), .ZN(n466) );
  and2 U571 ( .A1(n466), .A2(n536), .Z(n460) );
  or2 U572 ( .A1(n514), .A2(n466), .Z(n463) );
  inv1 U573 ( .I(n463), .ZN(n476) );
  or2 U574 ( .A1(n460), .A2(n476), .Z(n461) );
  and2 U575 ( .A1(n307), .A2(n461), .Z(d5) );
  or2 U576 ( .A1(m2), .A2(k2), .Z(n462) );
  and2 U577 ( .A1(n463), .A2(n462), .Z(n465) );
  or2 U578 ( .A1(c1), .A2(n275), .Z(n464) );
  or2 U579 ( .A1(n465), .A2(n464), .Z(n470) );
  or2 U580 ( .A1(c1), .A2(n466), .Z(n468) );
  inv1 U581 ( .I(n536), .ZN(n467) );
  or2 U582 ( .A1(n468), .A2(n467), .Z(n472) );
  or2 U583 ( .A1(n472), .A2(l2), .Z(n469) );
  and2 U584 ( .A1(n470), .A2(n469), .Z(n471) );
  inv1 U585 ( .I(n471), .ZN(e5) );
  inv1 U586 ( .I(n472), .ZN(n474) );
  and2 U587 ( .A1(n269), .A2(l2), .Z(n473) );
  and2 U588 ( .A1(n474), .A2(n473), .Z(n480) );
  and2 U589 ( .A1(m2), .A2(n307), .Z(n478) );
  or2 U590 ( .A1(n476), .A2(n275), .Z(n477) );
  and2 U591 ( .A1(n478), .A2(n477), .Z(n479) );
  or2 U592 ( .A1(n480), .A2(n479), .Z(f5) );
  and2 U594 ( .A1(n2), .A2(n307), .Z(n481) );
  and2 U595 ( .A1(n485), .A2(n481), .Z(n482) );
  or2 U596 ( .A1(n483), .A2(n482), .Z(g5) );
  and2 U597 ( .A1(n2), .A2(n528), .Z(n484) );
  and2 U598 ( .A1(n517), .A2(n484), .Z(n489) );
  and2 U599 ( .A1(n307), .A2(o2), .Z(n487) );
  and2 U601 ( .A1(n487), .A2(n486), .Z(n488) );
  or2 U602 ( .A1(n489), .A2(n488), .Z(h5) );
  inv1 U603 ( .I(p2), .ZN(n492) );
  inv1 U605 ( .I(n490), .ZN(n506) );
  and2 U606 ( .A1(n492), .A2(n506), .Z(n491) );
  and2 U607 ( .A1(n517), .A2(n491), .Z(n497) );
  and2 U608 ( .A1(n298), .A2(n506), .Z(n494) );
  or2 U609 ( .A1(c1), .A2(n492), .Z(n493) );
  or2 U610 ( .A1(n494), .A2(n493), .Z(n495) );
  inv1 U611 ( .I(n495), .ZN(n496) );
  or2 U612 ( .A1(n497), .A2(n496), .Z(i5) );
  and2 U613 ( .A1(p2), .A2(n506), .Z(n498) );
  inv1 U617 ( .I(n500), .ZN(n502) );
  inv1 U618 ( .I(q2), .ZN(n501) );
  or2 U619 ( .A1(n502), .A2(n501), .Z(n503) );
  and2 U621 ( .A1(q2), .A2(p2), .Z(n505) );
  and2 U622 ( .A1(n506), .A2(n505), .Z(n507) );
  inv1 U626 ( .I(n510), .ZN(n511) );
  or2 U627 ( .A1(n511), .A2(n520), .Z(n512) );
  and2 U628 ( .A1(n513), .A2(n512), .Z(k5) );
  and2 U629 ( .A1(n524), .A2(n536), .Z(n516) );
  or2 U630 ( .A1(n280), .A2(n537), .Z(n515) );
  and2 U631 ( .A1(n516), .A2(n515), .Z(n5) );
  inv1f U337 ( .I(m1), .ZN(n527) );
  inv1f U338 ( .I(n434), .ZN(n451) );
  inv1 U339 ( .I(n529), .ZN(n539) );
  inv1 U340 ( .I(n535), .ZN(n18) );
  and2 U341 ( .A1(a0), .A2(n451), .Z(n439) );
  and2 U343 ( .A1(c0), .A2(n451), .Z(n447) );
  or2f U344 ( .A1(n2), .A2(n528), .Z(n267) );
  or2 U345 ( .A1(n288), .A2(i0), .Z(n414) );
  inv1 U346 ( .I(n533), .ZN(n309) );
  or2 U349 ( .A1(n323), .A2(n314), .Z(n297) );
  inv1 U350 ( .I(m0), .ZN(n306) );
  inv1 U351 ( .I(g0), .ZN(n362) );
  inv1 U353 ( .I(n15), .ZN(n540) );
  inv1 U354 ( .I(n291), .ZN(n285) );
  inv1 U355 ( .I(n368), .ZN(n542) );
  or2 U357 ( .A1(n485), .A2(n522), .Z(n486) );
  and2 U358 ( .A1(u1), .A2(n544), .Z(n389) );
  or2 U359 ( .A1(n444), .A2(n443), .Z(n446) );
  and2 U361 ( .A1(n522), .A2(n517), .Z(n483) );
  and2 U362 ( .A1(n504), .A2(n503), .Z(j5) );
  or2f U363 ( .A1(n417), .A2(n416), .Z(n419) );
  and2 U365 ( .A1(v), .A2(n456), .Z(n416) );
  and2 U366 ( .A1(y), .A2(n456), .Z(n428) );
  and2 U367 ( .A1(w), .A2(n456), .Z(n420) );
  inv1 U368 ( .I(n2), .ZN(n525) );
  inv1 U369 ( .I(n2), .ZN(n522) );
  inv1f U371 ( .I(n533), .ZN(n526) );
  and2f U374 ( .A1(v1), .A2(n309), .Z(n390) );
  and2f U376 ( .A1(u1), .A2(n309), .Z(n385) );
  and2f U377 ( .A1(y1), .A2(n309), .Z(n402) );
  and2f U378 ( .A1(t1), .A2(n309), .Z(n381) );
  and2f U380 ( .A1(h2), .A2(n309), .Z(n445) );
  and2f U382 ( .A1(i2), .A2(n542), .Z(n449) );
  and2f U385 ( .A1(j2), .A2(n542), .Z(n454) );
  and2f U386 ( .A1(g2), .A2(n542), .Z(n441) );
  and2f U392 ( .A1(f2), .A2(n542), .Z(n437) );
  and2f U393 ( .A1(z1), .A2(n542), .Z(n406) );
  or2f U394 ( .A1(n347), .A2(m1), .Z(n348) );
  or2f U395 ( .A1(n322), .A2(n321), .Z(n323) );
  and2 U399 ( .A1(s), .A2(n302), .Z(n400) );
  and2 U404 ( .A1(p), .A2(n302), .Z(n388) );
  inv1f U407 ( .I(n364), .ZN(n302) );
  inv1f U410 ( .I(n361), .ZN(n408) );
  and2f U415 ( .A1(n284), .A2(i2), .Z(n453) );
  and2f U416 ( .A1(n284), .A2(g2), .Z(n444) );
  inv1f U427 ( .I(n270), .ZN(n544) );
  inv1 U428 ( .I(o2), .ZN(n528) );
  and2f U431 ( .A1(v2), .A2(g0), .Z(n271) );
  inv1f U432 ( .I(n270), .ZN(n301) );
  or2f U433 ( .A1(n241), .A2(n217), .Z(n238) );
  and2f U434 ( .A1(n284), .A2(t1), .Z(n384) );
  inv1 U439 ( .I(n361), .ZN(n284) );
  and2f U441 ( .A1(n408), .A2(w1), .Z(n397) );
  or2f U443 ( .A1(n421), .A2(n420), .Z(n423) );
  or2f U444 ( .A1(n429), .A2(n428), .Z(n431) );
  or2f U445 ( .A1(n453), .A2(n452), .Z(n455) );
  or2f U446 ( .A1(n265), .A2(n266), .Z(n529) );
  or2f U453 ( .A1(p2), .A2(n216), .Z(n265) );
  and2f U454 ( .A1(k), .A2(n387), .Z(n365) );
  or2f U455 ( .A1(n275), .A2(k2), .Z(n273) );
  inv1f U456 ( .I(l2), .ZN(n275) );
  and2f U458 ( .A1(z), .A2(n456), .Z(n435) );
  and2f U459 ( .A1(n169), .A2(n170), .Z(n165) );
  or2f U460 ( .A1(n389), .A2(n388), .Z(n391) );
  or2f U463 ( .A1(n380), .A2(n379), .Z(n382) );
  and2f U466 ( .A1(n285), .A2(s1), .Z(n380) );
  or2f U467 ( .A1(n393), .A2(n392), .Z(n395) );
  and2f U471 ( .A1(n285), .A2(v1), .Z(n393) );
  and2f U473 ( .A1(n285), .A2(a2), .Z(n417) );
  or2f U476 ( .A1(n425), .A2(n424), .Z(n427) );
  and2f U478 ( .A1(n285), .A2(c2), .Z(n425) );
  or2f U479 ( .A1(n440), .A2(n439), .Z(n442) );
  and2f U481 ( .A1(n285), .A2(f2), .Z(n440) );
  or2f U482 ( .A1(n448), .A2(n447), .Z(n450) );
  and2f U484 ( .A1(n285), .A2(h2), .Z(n448) );
  or2f U486 ( .A1(n376), .A2(n375), .Z(n378) );
  and2f U487 ( .A1(r1), .A2(n457), .Z(n376) );
  or2f U488 ( .A1(n405), .A2(n404), .Z(n407) );
  inv1f U489 ( .I(h0), .ZN(n531) );
  inv1 U491 ( .I(h0), .ZN(n530) );
  inv1f U493 ( .I(h0), .ZN(n350) );
  and2f U496 ( .A1(n354), .A2(n355), .Z(n532) );
  or2f U497 ( .A1(n292), .A2(n414), .Z(n415) );
  or2f U502 ( .A1(n367), .A2(n413), .Z(n533) );
  and2f U503 ( .A1(n279), .A2(n290), .Z(n413) );
  and2f U504 ( .A1(e1), .A2(n306), .Z(n534) );
  and2f U508 ( .A1(e1), .A2(n306), .Z(n288) );
  or2f U509 ( .A1(n320), .A2(n362), .Z(n324) );
  or2f U511 ( .A1(n362), .A2(n314), .Z(n342) );
  or2f U512 ( .A1(n362), .A2(i0), .Z(n294) );
  or2f U516 ( .A1(n265), .A2(n266), .Z(n535) );
  or2f U517 ( .A1(n523), .A2(n267), .Z(n266) );
  or2f U518 ( .A1(n276), .A2(n286), .Z(n335) );
  or2f U519 ( .A1(n530), .A2(g), .Z(n286) );
  or2 U520 ( .A1(n280), .A2(u2), .Z(n536) );
  or2f U521 ( .A1(n280), .A2(u2), .Z(n514) );
  and2f U525 ( .A1(n281), .A2(b), .Z(n280) );
  or2f U526 ( .A1(n314), .A2(n527), .Z(n315) );
  or2f U529 ( .A1(n527), .A2(n314), .Z(n293) );
  inv1f U531 ( .I(v2), .ZN(n314) );
  and2f U535 ( .A1(n271), .A2(m1), .Z(n354) );
  or2 U536 ( .A1(n339), .A2(k2), .Z(n537) );
  or2f U539 ( .A1(n339), .A2(k2), .Z(n272) );
  or2f U540 ( .A1(n275), .A2(n269), .Z(n339) );
  and2f U541 ( .A1(r), .A2(n302), .Z(n396) );
  and2f U542 ( .A1(l), .A2(n302), .Z(n371) );
  and2f U544 ( .A1(o), .A2(n302), .Z(n383) );
  or2f U546 ( .A1(n401), .A2(n400), .Z(n403) );
  inv1f U547 ( .I(n236), .ZN(n538) );
  or2f U548 ( .A1(n239), .A2(n238), .Z(n236) );
  inv1f U549 ( .I(n434), .ZN(n456) );
  inv1 U551 ( .I(n539), .ZN(n541) );
  and2f U552 ( .A1(m1), .A2(n530), .Z(n319) );
  and2f U553 ( .A1(n295), .A2(n296), .Z(n303) );
  or2f U554 ( .A1(n324), .A2(n297), .Z(n295) );
  or2f U556 ( .A1(n532), .A2(n414), .Z(n291) );
  and2f U557 ( .A1(n307), .A2(n499), .Z(n504) );
  or2f U558 ( .A1(n500), .A2(q2), .Z(n499) );
  and2f U559 ( .A1(n508), .A2(n498), .Z(n500) );
  and2f U561 ( .A1(n355), .A2(n279), .Z(n292) );
  and2f U563 ( .A1(n271), .A2(m1), .Z(n279) );
  or2f U564 ( .A1(n276), .A2(n327), .Z(n355) );
  or2f U570 ( .A1(n528), .A2(n522), .Z(n490) );
  and2f U593 ( .A1(p1), .A2(n301), .Z(n366) );
  and2f U600 ( .A1(z1), .A2(n457), .Z(n410) );
  and2f U604 ( .A1(e2), .A2(n457), .Z(n436) );
  and2f U614 ( .A1(q1), .A2(n301), .Z(n372) );
  or2f U615 ( .A1(n433), .A2(n432), .Z(n434) );
  inv1f U616 ( .I(n335), .ZN(n432) );
  and2f U620 ( .A1(b0), .A2(n451), .Z(n443) );
  or2f U623 ( .A1(n265), .A2(n266), .Z(n15) );
  or2f U624 ( .A1(n523), .A2(n525), .Z(n240) );
  and2f U625 ( .A1(u), .A2(n387), .Z(n409) );
  inv1f U632 ( .I(n364), .ZN(n387) );
  or2f U633 ( .A1(n299), .A2(n432), .Z(n364) );
  inv1f U634 ( .I(n533), .ZN(n543) );
  inv1f U635 ( .I(n368), .ZN(n308) );
  or2f U636 ( .A1(n367), .A2(n413), .Z(n368) );
  and2f U637 ( .A1(n307), .A2(n509), .Z(n513) );
  or2f U638 ( .A1(n510), .A2(r2), .Z(n509) );
  and2f U639 ( .A1(n508), .A2(n507), .Z(n510) );
  or2f U640 ( .A1(n274), .A2(n340), .Z(n508) );
  inv1f U641 ( .I(n298), .ZN(n485) );
  or2f U642 ( .A1(n343), .A2(n340), .Z(n298) );
  inv1f U643 ( .I(n341), .ZN(n517) );
  or2f U644 ( .A1(n485), .A2(c1), .Z(n341) );
  or2f U645 ( .A1(n300), .A2(n414), .Z(n361) );
  and2f U646 ( .A1(n354), .A2(n355), .Z(n300) );
  or2f U647 ( .A1(n292), .A2(n414), .Z(n270) );
  inv1f U648 ( .I(n415), .ZN(n457) );
endmodule

