
module C1908_iscas ( g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, 
        p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, f1, e1, d1, c1, b1, a1, 
        z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, 
        h0 );
  input g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m,
         l, k, j, i, h, g, f, e, d, c, b, a;
  output f1, e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0,
         o0, n0, m0, l0, k0, j0, i0, h0;
  wire   n256, n366, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n503, n504, n505, n506, n507, n508, n509, n511, n512, n513,
         n514, n516, n517, n518, n519, n520, n521, n522, n523, n524, n526,
         n527, n528, n529, n530, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n567, n568, n569, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n587, n588,
         n589, n590, n591, n592, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n633, n634, n635, n636, n637,
         n638, n639, n640, n642, n643, n645, n646, n647, n648, n649, n650,
         n651, n652, n654, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n730, n731, n732,
         n734, n735, n736, n737, n738, n739, n741, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1013,
         n1014, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1110, n1111, n1112, n1113, n1114, n1115, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275;

  or2 U341 ( .A1(n256), .A2(n1275), .Z(n366) );
  and2 U345 ( .A1(w), .A2(x), .Z(n256) );
  and2 U493 ( .A1(n597), .A2(n598), .Z(n468) );
  or2 U494 ( .A1(n995), .A2(n996), .Z(n469) );
  and2 U495 ( .A1(n627), .A2(n628), .Z(n470) );
  or2 U497 ( .A1(n493), .A2(n1019), .Z(n471) );
  or2 U498 ( .A1(n519), .A2(n518), .Z(n472) );
  and2 U499 ( .A1(j), .A2(n1014), .Z(n473) );
  or2 U511 ( .A1(n1189), .A2(n1190), .Z(c1) );
  or2 U514 ( .A1(n1086), .A2(n622), .Z(n482) );
  or2 U517 ( .A1(n507), .A2(n485), .Z(n602) );
  or2 U520 ( .A1(n1230), .A2(n768), .Z(n487) );
  or2 U523 ( .A1(n1036), .A2(n1038), .Z(n489) );
  and2 U525 ( .A1(n678), .A2(o), .Z(n491) );
  and2 U528 ( .A1(n909), .A2(n496), .Z(n494) );
  and2 U530 ( .A1(n812), .A2(n810), .Z(n495) );
  and2 U531 ( .A1(n808), .A2(n812), .Z(n496) );
  or2 U533 ( .A1(n499), .A2(n500), .Z(n498) );
  inv1 U534 ( .I(n627), .ZN(n499) );
  inv1 U535 ( .I(n628), .ZN(n500) );
  or2 U536 ( .A1(n1085), .A2(n490), .Z(n501) );
  inv1 U540 ( .I(n504), .ZN(n674) );
  or2 U541 ( .A1(n1173), .A2(n841), .Z(n505) );
  inv1 U544 ( .I(n776), .ZN(n507) );
  or2 U552 ( .A1(n981), .A2(n552), .Z(n514) );
  or2 U554 ( .A1(n791), .A2(n790), .Z(n516) );
  inv1 U557 ( .I(n544), .ZN(n519) );
  or2 U559 ( .A1(n804), .A2(n968), .Z(n521) );
  inv1 U572 ( .I(n1076), .ZN(n533) );
  and2 U575 ( .A1(n645), .A2(n898), .Z(n537) );
  inv1 U579 ( .I(n539), .ZN(n1245) );
  and2 U581 ( .A1(n761), .A2(n1159), .Z(n541) );
  inv1 U583 ( .I(n542), .ZN(n1164) );
  inv1 U584 ( .I(n541), .ZN(n543) );
  inv1 U587 ( .I(n545), .ZN(n1076) );
  or2 U590 ( .A1(n815), .A2(e0), .Z(n548) );
  or2 U593 ( .A1(n1239), .A2(n968), .Z(n550) );
  or2 U600 ( .A1(e0), .A2(n940), .Z(n555) );
  inv1 U603 ( .I(n558), .ZN(n1123) );
  or2 U605 ( .A1(n1121), .A2(n551), .Z(n560) );
  or2 U607 ( .A1(n807), .A2(a), .Z(n562) );
  and2 U609 ( .A1(n816), .A2(n691), .Z(n564) );
  and2 U612 ( .A1(n595), .A2(p), .Z(n567) );
  and2 U613 ( .A1(n), .A2(n767), .Z(n568) );
  and2 U614 ( .A1(p), .A2(n595), .Z(n569) );
  and2 U616 ( .A1(n887), .A2(n573), .Z(n571) );
  or2 U617 ( .A1(n571), .A2(n572), .Z(n650) );
  or2 U623 ( .A1(n578), .A2(k), .Z(n577) );
  inv1 U624 ( .I(n914), .ZN(n578) );
  inv1 U626 ( .I(n666), .ZN(n580) );
  or2 U627 ( .A1(n745), .A2(n886), .Z(n581) );
  or2 U628 ( .A1(n621), .A2(n583), .Z(n582) );
  inv1 U630 ( .I(n866), .ZN(n583) );
  or2 U633 ( .A1(n756), .A2(n589), .Z(n587) );
  or2 U635 ( .A1(n777), .A2(n583), .Z(n588) );
  and2 U637 ( .A1(o), .A2(n1007), .Z(n590) );
  and2 U640 ( .A1(j), .A2(n764), .Z(n592) );
  and2 U642 ( .A1(n595), .A2(p), .Z(n594) );
  and2 U644 ( .A1(n887), .A2(n886), .Z(n596) );
  or2 U645 ( .A1(n599), .A2(n943), .Z(n597) );
  and2 U646 ( .A1(n597), .A2(n598), .Z(n952) );
  or2 U647 ( .A1(e0), .A2(n724), .Z(n598) );
  or2 U648 ( .A1(n995), .A2(n996), .Z(n600) );
  or2 U649 ( .A1(n1011), .A2(n530), .Z(n601) );
  inv1 U651 ( .I(n622), .ZN(n604) );
  inv1 U654 ( .I(n574), .ZN(n1008) );
  or2 U657 ( .A1(n1266), .A2(n762), .Z(n609) );
  and2 U658 ( .A1(n624), .A2(n611), .Z(n610) );
  inv1 U659 ( .I(n609), .ZN(n611) );
  or2 U660 ( .A1(n563), .A2(n1085), .Z(n612) );
  inv1 U662 ( .I(n613), .ZN(n937) );
  and2 U669 ( .A1(n732), .A2(n968), .Z(n619) );
  and2 U670 ( .A1(n787), .A2(n767), .Z(n620) );
  or2 U671 ( .A1(n756), .A2(n865), .Z(n621) );
  or2 U673 ( .A1(n596), .A2(n623), .Z(n645) );
  or2 U674 ( .A1(n889), .A2(n737), .Z(n623) );
  or2 U688 ( .A1(n757), .A2(n1038), .Z(n637) );
  or2 U690 ( .A1(n1084), .A2(n648), .Z(n638) );
  inv1 U691 ( .I(n969), .ZN(n639) );
  and2 U692 ( .A1(n867), .A2(n583), .Z(n640) );
  inv1 U694 ( .I(n976), .ZN(n642) );
  inv1 U696 ( .I(c), .ZN(n643) );
  inv1 U697 ( .I(n645), .ZN(n670) );
  or2 U699 ( .A1(n968), .A2(n805), .Z(n647) );
  inv1 U701 ( .I(n600), .ZN(n649) );
  or2 U703 ( .A1(n1040), .A2(n575), .Z(n652) );
  and2 U711 ( .A1(n767), .A2(n1234), .Z(n658) );
  or2 U713 ( .A1(n919), .A2(n660), .Z(n926) );
  inv1 U716 ( .I(n661), .ZN(n791) );
  inv1 U718 ( .I(p), .ZN(n663) );
  and2 U721 ( .A1(n667), .A2(n1185), .Z(n666) );
  inv1 U722 ( .I(n1183), .ZN(n667) );
  and2 U726 ( .A1(n694), .A2(m), .Z(n675) );
  and2 U729 ( .A1(n678), .A2(o), .Z(n677) );
  inv1 U730 ( .I(j), .ZN(n678) );
  and2 U734 ( .A1(n722), .A2(l), .Z(n681) );
  or2 U738 ( .A1(n639), .A2(n1130), .Z(n685) );
  or2 U739 ( .A1(n734), .A2(b), .Z(n686) );
  and2 U741 ( .A1(n734), .A2(b), .Z(n688) );
  inv1 U742 ( .I(n936), .ZN(n689) );
  and2 U743 ( .A1(n691), .A2(n816), .Z(n690) );
  inv1 U744 ( .I(n1138), .ZN(n691) );
  inv1 U745 ( .I(n486), .ZN(n984) );
  inv1 U749 ( .I(l), .ZN(n694) );
  or2 U753 ( .A1(n786), .A2(n767), .Z(n698) );
  or2 U757 ( .A1(n815), .A2(e0), .Z(n701) );
  or2 U758 ( .A1(n810), .A2(n812), .Z(n702) );
  inv1 U759 ( .I(f), .ZN(n703) );
  or2 U760 ( .A1(n702), .A2(n809), .Z(n704) );
  inv1 U763 ( .I(n705), .ZN(n928) );
  or2 U765 ( .A1(n791), .A2(n708), .Z(n707) );
  or2 U767 ( .A1(n633), .A2(n657), .Z(n708) );
  and2 U769 ( .A1(p), .A2(n711), .Z(n710) );
  inv1 U770 ( .I(n), .ZN(n711) );
  inv1 U774 ( .I(n714), .ZN(n808) );
  inv1 U778 ( .I(n1139), .ZN(n717) );
  inv1 U781 ( .I(n1167), .ZN(n719) );
  inv1 U783 ( .I(n720), .ZN(n1181) );
  inv1 U784 ( .I(n1175), .ZN(n721) );
  inv1 U785 ( .I(m), .ZN(n722) );
  and2 U786 ( .A1(n950), .A2(n724), .Z(n723) );
  inv1 U787 ( .I(n951), .ZN(n724) );
  and2 U792 ( .A1(b), .A2(n859), .Z(n728) );
  or2 U794 ( .A1(n695), .A2(n662), .Z(n730) );
  inv1 U795 ( .I(n730), .ZN(n862) );
  inv1 U796 ( .I(p), .ZN(n731) );
  or2 U797 ( .A1(n915), .A2(n682), .Z(n732) );
  inv1 U800 ( .I(c), .ZN(n734) );
  or2 U801 ( .A1(n569), .A2(n860), .Z(n735) );
  and2 U802 ( .A1(n753), .A2(n737), .Z(n736) );
  or2 U804 ( .A1(n1025), .A2(n1024), .Z(n738) );
  inv1 U805 ( .I(n738), .ZN(n739) );
  or2 U811 ( .A1(n581), .A2(n746), .Z(n744) );
  and2 U812 ( .A1(n879), .A2(n747), .Z(n745) );
  or2 U813 ( .A1(n745), .A2(n746), .Z(n884) );
  and2 U814 ( .A1(n881), .A2(n997), .Z(n746) );
  and2 U815 ( .A1(i), .A2(n997), .Z(n747) );
  or2 U819 ( .A1(n1052), .A2(n1087), .Z(n749) );
  or2 U822 ( .A1(e0), .A2(n1165), .Z(n751) );
  inv1 U831 ( .I(n1141), .ZN(n760) );
  inv1 U832 ( .I(n1158), .ZN(n761) );
  inv1 U833 ( .I(n579), .ZN(n1190) );
  inv1 U834 ( .I(n1268), .ZN(n762) );
  or2 U838 ( .A1(n698), .A2(n590), .Z(n766) );
  inv1 U840 ( .I(p), .ZN(n767) );
  or2 U846 ( .A1(n774), .A2(n728), .Z(n773) );
  inv1 U850 ( .I(n776), .ZN(n872) );
  inv1 U852 ( .I(n778), .ZN(n1084) );
  or2 U853 ( .A1(n507), .A2(n687), .Z(n779) );
  or2 U855 ( .A1(n1040), .A2(n575), .Z(n781) );
  inv1 U857 ( .I(n1137), .ZN(n783) );
  or2 U858 ( .A1(n757), .A2(n1057), .Z(n784) );
  inv1 U859 ( .I(e0), .ZN(n1275) );
  or2 U860 ( .A1(e0), .A2(x), .Z(n785) );
  inv1 U861 ( .I(n785), .ZN(n962) );
  inv1 U862 ( .I(q), .ZN(n904) );
  or2 U863 ( .A1(n962), .A2(n904), .Z(n1138) );
  inv1 U864 ( .I(o), .ZN(n1014) );
  and2 U868 ( .A1(n524), .A2(n767), .Z(n788) );
  inv1 U870 ( .I(i), .ZN(n1234) );
  inv1 U871 ( .I(u), .ZN(n792) );
  or2 U872 ( .A1(g0), .A2(n792), .Z(n1142) );
  inv1 U873 ( .I(n1142), .ZN(n1140) );
  inv1 U875 ( .I(n516), .ZN(n1145) );
  inv1 U876 ( .I(d), .ZN(n997) );
  and2 U877 ( .A1(h), .A2(n997), .Z(n796) );
  and2 U878 ( .A1(n528), .A2(d), .Z(n795) );
  or2 U879 ( .A1(n796), .A2(n795), .Z(n811) );
  or2 U881 ( .A1(n1041), .A2(f), .Z(n800) );
  inv1 U882 ( .I(f), .ZN(n1032) );
  or2 U883 ( .A1(g), .A2(n703), .Z(n799) );
  and2 U884 ( .A1(n800), .A2(n799), .Z(n797) );
  or2 U885 ( .A1(n797), .A2(e), .Z(n798) );
  inv1 U886 ( .I(n798), .ZN(n803) );
  inv1 U890 ( .I(a), .ZN(n968) );
  inv1 U891 ( .I(b), .ZN(n975) );
  inv1 U892 ( .I(c), .ZN(n983) );
  or2 U893 ( .A1(n643), .A2(b), .Z(n806) );
  inv1 U894 ( .I(n806), .ZN(n804) );
  or2 U895 ( .A1(n688), .A2(n804), .Z(n805) );
  or2 U897 ( .A1(n807), .A2(a), .Z(n934) );
  and2 U900 ( .A1(n909), .A2(n808), .Z(n809) );
  inv1 U901 ( .I(n811), .ZN(n812) );
  inv1 U905 ( .I(l), .ZN(n1066) );
  and2 U906 ( .A1(o), .A2(n1066), .Z(n818) );
  and2 U907 ( .A1(n764), .A2(l), .Z(n817) );
  or2 U908 ( .A1(n818), .A2(n817), .Z(n822) );
  and2 U909 ( .A1(n528), .A2(j), .Z(n820) );
  or2 U911 ( .A1(n820), .A2(n819), .Z(n823) );
  inv1 U912 ( .I(n823), .ZN(n821) );
  and2 U913 ( .A1(n822), .A2(n821), .Z(n826) );
  inv1 U914 ( .I(n822), .ZN(n824) );
  and2 U915 ( .A1(n824), .A2(n823), .Z(n825) );
  and2 U917 ( .A1(f), .A2(n983), .Z(n828) );
  inv1 U922 ( .I(s), .ZN(n877) );
  inv1 U924 ( .I(n831), .ZN(n829) );
  and2 U927 ( .A1(n832), .A2(n831), .Z(n833) );
  or2 U928 ( .A1(n834), .A2(n833), .Z(n837) );
  inv1 U929 ( .I(n837), .ZN(n835) );
  inv1 U931 ( .I(n836), .ZN(n838) );
  or2 U933 ( .A1(n840), .A2(n839), .Z(n1176) );
  inv1 U935 ( .I(b0), .ZN(n1173) );
  and2 U936 ( .A1(n1173), .A2(n841), .Z(n842) );
  inv1 U938 ( .I(k), .ZN(n1060) );
  and2 U939 ( .A1(o), .A2(n1060), .Z(n845) );
  and2 U940 ( .A1(n764), .A2(k), .Z(n844) );
  or2 U941 ( .A1(n845), .A2(n844), .Z(n849) );
  inv1 U942 ( .I(e), .ZN(n1026) );
  and2 U943 ( .A1(h), .A2(n1026), .Z(n847) );
  or2 U945 ( .A1(n847), .A2(n846), .Z(n850) );
  inv1 U946 ( .I(n850), .ZN(n848) );
  and2 U947 ( .A1(n849), .A2(n848), .Z(n853) );
  inv1 U948 ( .I(n849), .ZN(n851) );
  and2 U949 ( .A1(n851), .A2(n850), .Z(n852) );
  or2 U951 ( .A1(g0), .A2(x), .Z(n905) );
  inv1 U952 ( .I(r), .ZN(n961) );
  or2 U953 ( .A1(n905), .A2(n961), .Z(n866) );
  and2 U955 ( .A1(n), .A2(n731), .Z(n854) );
  or2 U956 ( .A1(n567), .A2(n854), .Z(n856) );
  inv1 U957 ( .I(n856), .ZN(n855) );
  and2 U962 ( .A1(n731), .A2(n), .Z(n860) );
  and2 U968 ( .A1(n870), .A2(n777), .Z(n871) );
  inv1 U969 ( .I(a0), .ZN(n1165) );
  or2 U974 ( .A1(n769), .A2(n616), .Z(n932) );
  or2 U975 ( .A1(e0), .A2(n875), .Z(n876) );
  inv1 U976 ( .I(n876), .ZN(n958) );
  or2 U977 ( .A1(n958), .A2(n877), .Z(n1182) );
  and2 U978 ( .A1(n1275), .A2(n1182), .Z(n898) );
  or2 U984 ( .A1(n882), .A2(n881), .Z(n883) );
  or2 U985 ( .A1(n671), .A2(n884), .Z(n887) );
  inv1 U986 ( .I(t), .ZN(n957) );
  or2 U987 ( .A1(n885), .A2(n957), .Z(n888) );
  inv1 U988 ( .I(n888), .ZN(n886) );
  and2 U989 ( .A1(n887), .A2(n886), .Z(n890) );
  inv1 U991 ( .I(m), .ZN(n1071) );
  and2 U992 ( .A1(j), .A2(n1071), .Z(n891) );
  or2 U993 ( .A1(n892), .A2(n891), .Z(n893) );
  and2 U994 ( .A1(n1041), .A2(n893), .Z(n896) );
  inv1 U995 ( .I(n893), .ZN(n894) );
  and2 U996 ( .A1(g), .A2(n894), .Z(n895) );
  or2 U997 ( .A1(n896), .A2(n895), .Z(n897) );
  or2 U998 ( .A1(n670), .A2(n736), .Z(n1184) );
  inv1 U999 ( .I(n1184), .ZN(n1186) );
  inv1 U1001 ( .I(n1182), .ZN(n901) );
  or2 U1002 ( .A1(n650), .A2(e0), .Z(n899) );
  or2 U1005 ( .A1(n905), .A2(n904), .Z(n908) );
  inv1 U1006 ( .I(n908), .ZN(n906) );
  and2 U1007 ( .A1(n713), .A2(n906), .Z(n911) );
  and2 U1010 ( .A1(n694), .A2(m), .Z(n913) );
  and2 U1011 ( .A1(n722), .A2(l), .Z(n912) );
  inv1 U1016 ( .I(n1239), .ZN(n1241) );
  inv1 U1021 ( .I(z), .ZN(n1265) );
  or2 U1022 ( .A1(e0), .A2(n1265), .Z(n924) );
  inv1 U1024 ( .I(n925), .ZN(n972) );
  inv1 U1032 ( .I(v), .ZN(n939) );
  or2 U1033 ( .A1(g0), .A2(n939), .Z(n942) );
  inv1 U1034 ( .I(n942), .ZN(n940) );
  or2 U1035 ( .A1(n943), .A2(n741), .Z(n950) );
  and2 U1036 ( .A1(n997), .A2(n), .Z(n945) );
  and2 U1037 ( .A1(d), .A2(n595), .Z(n944) );
  or2 U1038 ( .A1(n945), .A2(n944), .Z(n946) );
  and2 U1039 ( .A1(n946), .A2(n584), .Z(n949) );
  inv1 U1040 ( .I(n946), .ZN(n947) );
  and2 U1041 ( .A1(n947), .A2(n483), .Z(n948) );
  or2 U1042 ( .A1(n949), .A2(n948), .Z(n951) );
  inv1 U1044 ( .I(y), .ZN(n1157) );
  or2 U1049 ( .A1(n958), .A2(n957), .Z(n959) );
  inv1 U1050 ( .I(n959), .ZN(n1038) );
  or2 U1052 ( .A1(n962), .A2(n961), .Z(n1082) );
  inv1 U1053 ( .I(n1082), .ZN(n1087) );
  inv1 U1054 ( .I(f0), .ZN(n963) );
  or2 U1055 ( .A1(g0), .A2(n963), .Z(n1002) );
  or2 U1056 ( .A1(n1002), .A2(n256), .Z(n966) );
  inv1 U1057 ( .I(g0), .ZN(n1227) );
  or2 U1058 ( .A1(n1227), .A2(c0), .Z(n964) );
  or2 U1059 ( .A1(n964), .A2(n366), .Z(n965) );
  and2 U1060 ( .A1(n966), .A2(n965), .Z(n967) );
  or2 U1061 ( .A1(n1087), .A2(n967), .Z(n1036) );
  or2 U1065 ( .A1(n639), .A2(a), .Z(n971) );
  or2 U1066 ( .A1(n969), .A2(n968), .Z(n970) );
  and2 U1067 ( .A1(n971), .A2(n970), .Z(h0) );
  or2 U1069 ( .A1(n659), .A2(n1085), .Z(n1018) );
  or2 U1070 ( .A1(n973), .A2(n972), .Z(n1094) );
  inv1 U1074 ( .I(n976), .ZN(n1130) );
  or2 U1075 ( .A1(n1130), .A2(b), .Z(n978) );
  or2 U1076 ( .A1(n976), .A2(n975), .Z(n977) );
  and2 U1077 ( .A1(n978), .A2(n977), .Z(i0) );
  or2 U1078 ( .A1(n1037), .A2(n1084), .Z(n980) );
  or2 U1079 ( .A1(n517), .A2(n980), .Z(n982) );
  inv1 U1080 ( .I(n984), .ZN(n1199) );
  or2 U1081 ( .A1(n1199), .A2(c), .Z(n986) );
  or2 U1082 ( .A1(n984), .A2(n734), .Z(n985) );
  and2 U1083 ( .A1(n986), .A2(n985), .Z(j0) );
  or2 U1086 ( .A1(n664), .A2(n1036), .Z(n993) );
  or2 U1087 ( .A1(n755), .A2(n553), .Z(n991) );
  or2 U1088 ( .A1(n989), .A2(n553), .Z(n990) );
  or2 U1093 ( .A1(n1196), .A2(d), .Z(n999) );
  or2 U1094 ( .A1(n469), .A2(n997), .Z(n998) );
  and2 U1095 ( .A1(n999), .A2(n998), .Z(k0) );
  or2 U1096 ( .A1(n1275), .A2(n1227), .Z(n1000) );
  or2 U1097 ( .A1(n1000), .A2(d0), .Z(n1001) );
  and2 U1098 ( .A1(n1002), .A2(n1001), .Z(n1003) );
  or2 U1099 ( .A1(n1003), .A2(n256), .Z(n1052) );
  or2 U1100 ( .A1(n1052), .A2(n1087), .Z(n1057) );
  or2 U1101 ( .A1(n659), .A2(n1057), .Z(n1004) );
  or2 U1104 ( .A1(n574), .A2(j), .Z(n1010) );
  or2 U1105 ( .A1(n1008), .A2(n1007), .Z(n1009) );
  and2 U1106 ( .A1(n1010), .A2(n1009), .Z(l0) );
  or2 U1107 ( .A1(n530), .A2(n1011), .Z(n1045) );
  or2 U1108 ( .A1(n1045), .A2(n769), .Z(n1013) );
  inv1 U1110 ( .I(n477), .ZN(n1220) );
  or2 U1111 ( .A1(n1220), .A2(o), .Z(n1017) );
  or2 U1112 ( .A1(n477), .A2(n764), .Z(n1016) );
  and2 U1113 ( .A1(n1017), .A2(n1016), .Z(m0) );
  or2 U1114 ( .A1(n731), .A2(n1020), .Z(n1022) );
  or2 U1116 ( .A1(n696), .A2(p), .Z(n1021) );
  and2 U1117 ( .A1(n1022), .A2(n1021), .Z(n0) );
  or2 U1119 ( .A1(n679), .A2(n489), .Z(n1031) );
  or2 U1120 ( .A1(n1031), .A2(n1085), .Z(n1025) );
  or2 U1122 ( .A1(n1024), .A2(n612), .Z(n1027) );
  inv1 U1123 ( .I(n1027), .ZN(n1200) );
  or2 U1124 ( .A1(n1200), .A2(e), .Z(n1029) );
  or2 U1125 ( .A1(n1027), .A2(n1026), .Z(n1028) );
  and2 U1126 ( .A1(n1029), .A2(n1028), .Z(o0) );
  or2 U1129 ( .A1(n646), .A2(f), .Z(n1035) );
  or2 U1130 ( .A1(n513), .A2(n1032), .Z(n1034) );
  and2 U1131 ( .A1(n1035), .A2(n1034), .Z(p0) );
  or2 U1136 ( .A1(n634), .A2(n652), .Z(n1042) );
  inv1 U1137 ( .I(n1042), .ZN(n1132) );
  or2 U1138 ( .A1(n1132), .A2(g), .Z(n1044) );
  or2 U1139 ( .A1(n1042), .A2(n1041), .Z(n1043) );
  and2 U1140 ( .A1(n1044), .A2(n1043), .Z(q0) );
  or2 U1144 ( .A1(n1205), .A2(h), .Z(n1049) );
  or2 U1145 ( .A1(n1047), .A2(n528), .Z(n1048) );
  and2 U1146 ( .A1(n1049), .A2(n1048), .Z(r0) );
  or2 U1148 ( .A1(n1080), .A2(n1052), .Z(n1053) );
  or2 U1151 ( .A1(n1126), .A2(i), .Z(n1056) );
  or2 U1152 ( .A1(n1054), .A2(n1234), .Z(n1055) );
  and2 U1153 ( .A1(n1056), .A2(n1055), .Z(s0) );
  or2 U1154 ( .A1(n960), .A2(n784), .Z(n1058) );
  or2 U1155 ( .A1(n1245), .A2(n552), .Z(n1064) );
  or2 U1156 ( .A1(n1064), .A2(n1085), .Z(n1061) );
  inv1 U1157 ( .I(n1061), .ZN(n1059) );
  or2 U1158 ( .A1(n1059), .A2(k), .Z(n1063) );
  or2 U1159 ( .A1(n1061), .A2(n1060), .Z(n1062) );
  and2 U1160 ( .A1(n1063), .A2(n1062), .Z(t0) );
  or2 U1161 ( .A1(n1064), .A2(n604), .Z(n1067) );
  inv1 U1162 ( .I(n1067), .ZN(n1065) );
  or2 U1163 ( .A1(n1065), .A2(l), .Z(n1069) );
  or2 U1164 ( .A1(n1067), .A2(n1066), .Z(n1068) );
  and2 U1165 ( .A1(n1069), .A2(n1068), .Z(u0) );
  or2 U1166 ( .A1(n1245), .A2(n652), .Z(n1072) );
  inv1 U1167 ( .I(n1072), .ZN(n1070) );
  or2 U1168 ( .A1(n1070), .A2(m), .Z(n1074) );
  or2 U1169 ( .A1(n1072), .A2(n1071), .Z(n1073) );
  and2 U1170 ( .A1(n1074), .A2(n1073), .Z(v0) );
  or2 U1171 ( .A1(n533), .A2(n), .Z(n1078) );
  or2 U1172 ( .A1(n1076), .A2(n595), .Z(n1077) );
  and2 U1173 ( .A1(n1078), .A2(n1077), .Z(w0) );
  inv1 U1174 ( .I(n256), .ZN(n1079) );
  and2 U1175 ( .A1(n1079), .A2(f0), .Z(n1108) );
  inv1 U1177 ( .I(n1080), .ZN(n1112) );
  and2 U1178 ( .A1(n561), .A2(n1112), .Z(n1092) );
  inv1 U1179 ( .I(n616), .ZN(n1110) );
  or2 U1180 ( .A1(n768), .A2(n1082), .Z(n1083) );
  and2 U1181 ( .A1(n1110), .A2(n1083), .Z(n1090) );
  or2 U1184 ( .A1(n1233), .A2(n1087), .Z(n1088) );
  inv1 U1185 ( .I(n1088), .ZN(n1111) );
  and2 U1186 ( .A1(n482), .A2(n1111), .Z(n1089) );
  or2 U1187 ( .A1(n1090), .A2(n1089), .Z(n1091) );
  and2 U1188 ( .A1(n1092), .A2(n1091), .Z(n1106) );
  and2 U1189 ( .A1(n1110), .A2(n1111), .Z(n1104) );
  inv1 U1190 ( .I(n551), .ZN(n1093) );
  or2 U1191 ( .A1(n575), .A2(n1093), .Z(n1095) );
  and2 U1192 ( .A1(n1112), .A2(n1095), .Z(n1102) );
  or2 U1194 ( .A1(n1097), .A2(n648), .Z(n1099) );
  or2 U1195 ( .A1(n1099), .A2(n757), .Z(n1100) );
  or2 U1197 ( .A1(n1102), .A2(n1101), .Z(n1103) );
  and2 U1198 ( .A1(n1104), .A2(n1103), .Z(n1105) );
  and2 U1200 ( .A1(n1108), .A2(n1107), .Z(n1136) );
  and2 U1201 ( .A1(n1110), .A2(n561), .Z(n1114) );
  and2 U1202 ( .A1(n1112), .A2(n1111), .Z(n1113) );
  and2 U1203 ( .A1(n1114), .A2(n1113), .Z(n1115) );
  or2 U1204 ( .A1(n1115), .A2(g0), .Z(n1134) );
  inv1 U1209 ( .I(n652), .ZN(n1246) );
  inv1 U1210 ( .I(n493), .ZN(n1122) );
  or2 U1221 ( .A1(n1136), .A2(n1135), .Z(x0) );
  or2 U1223 ( .A1(n1275), .A2(n1138), .Z(n1139) );
  and2 U1224 ( .A1(n1140), .A2(n760), .Z(n1144) );
  and2 U1225 ( .A1(n1142), .A2(n1141), .Z(n1143) );
  or2 U1226 ( .A1(n1144), .A2(n1143), .Z(n1146) );
  and2 U1227 ( .A1(n1145), .A2(n1146), .Z(n1149) );
  inv1 U1228 ( .I(n1146), .ZN(n1147) );
  and2 U1229 ( .A1(n516), .A2(n1147), .Z(n1148) );
  or2 U1230 ( .A1(n1149), .A2(n1148), .Z(n1151) );
  or2 U1231 ( .A1(n1227), .A2(f0), .Z(n1270) );
  and2 U1232 ( .A1(n1151), .A2(n1270), .Z(n1150) );
  inv1 U1234 ( .I(n1151), .ZN(n1152) );
  and2 U1235 ( .A1(n1152), .A2(n1270), .Z(n1154) );
  or2 U1237 ( .A1(n1155), .A2(n1156), .Z(y0) );
  or2 U1238 ( .A1(n1157), .A2(n1275), .Z(n1158) );
  or2 U1239 ( .A1(n668), .A2(n723), .Z(n1160) );
  and2 U1240 ( .A1(n1270), .A2(n1160), .Z(n1159) );
  inv1 U1241 ( .I(n1160), .ZN(n1161) );
  and2 U1242 ( .A1(n1270), .A2(n1161), .Z(n1162) );
  or2 U1244 ( .A1(n1163), .A2(n1164), .Z(z0) );
  or2 U1245 ( .A1(n1165), .A2(n1275), .Z(n1166) );
  and2 U1247 ( .A1(n779), .A2(n1270), .Z(n1167) );
  inv1 U1248 ( .I(n779), .ZN(n1168) );
  and2 U1249 ( .A1(n1168), .A2(n1270), .Z(n1170) );
  or2 U1252 ( .A1(n1173), .A2(n1275), .Z(n1174) );
  and2 U1254 ( .A1(n1176), .A2(n1270), .Z(n1175) );
  inv1 U1255 ( .I(n1176), .ZN(n1177) );
  and2 U1256 ( .A1(n1177), .A2(n1270), .Z(n1179) );
  or2 U1258 ( .A1(n1181), .A2(n1180), .Z(b1) );
  or2 U1259 ( .A1(n1275), .A2(n1182), .Z(n1183) );
  and2 U1261 ( .A1(n1184), .A2(n1270), .Z(n1185) );
  and2 U1262 ( .A1(n1186), .A2(n1270), .Z(n1188) );
  and2 U1264 ( .A1(u), .A2(c0), .Z(n1191) );
  or2 U1265 ( .A1(n1191), .A2(n1227), .Z(n1212) );
  inv1 U1266 ( .I(c0), .ZN(n1192) );
  or2 U1267 ( .A1(n1227), .A2(n1192), .Z(n1195) );
  or2 U1270 ( .A1(n1196), .A2(n760), .Z(n1197) );
  or2 U1271 ( .A1(n1198), .A2(n1197), .Z(n1202) );
  or2 U1272 ( .A1(n1200), .A2(n1199), .Z(n1201) );
  inv1 U1274 ( .I(n634), .ZN(n1204) );
  and2 U1275 ( .A1(n1246), .A2(n1204), .Z(n1206) );
  or2 U1276 ( .A1(n1205), .A2(n1206), .Z(n1208) );
  or2 U1277 ( .A1(n1208), .A2(n685), .Z(n1209) );
  or2 U1278 ( .A1(n1212), .A2(n626), .Z(n1218) );
  inv1 U1280 ( .I(n1212), .ZN(n1213) );
  or2 U1281 ( .A1(n1214), .A2(n1213), .Z(n1216) );
  inv1 U1282 ( .I(n626), .ZN(n1215) );
  and2 U1284 ( .A1(n1217), .A2(n1218), .Z(d1) );
  and2 U1285 ( .A1(d0), .A2(v), .Z(n1219) );
  or2 U1286 ( .A1(n1219), .A2(n1227), .Z(n1256) );
  or2 U1289 ( .A1(n763), .A2(n696), .Z(n1224) );
  or2 U1290 ( .A1(n1225), .A2(n1224), .Z(n1229) );
  inv1 U1291 ( .I(d0), .ZN(n1226) );
  or2 U1292 ( .A1(n1227), .A2(n1226), .Z(n1228) );
  inv1 U1295 ( .I(n1051), .ZN(n1247) );
  and2 U1298 ( .A1(n1234), .A2(n), .Z(n1237) );
  and2 U1299 ( .A1(i), .A2(n595), .Z(n1236) );
  or2 U1300 ( .A1(n1237), .A2(n1236), .Z(n1240) );
  inv1 U1301 ( .I(n1240), .ZN(n1238) );
  and2 U1302 ( .A1(n1239), .A2(n1238), .Z(n1243) );
  and2 U1303 ( .A1(n1241), .A2(n1240), .Z(n1242) );
  or2 U1304 ( .A1(n1243), .A2(n1242), .Z(n1257) );
  or2 U1305 ( .A1(n1244), .A2(n1257), .Z(n1252) );
  and2 U1307 ( .A1(n1246), .A2(n539), .Z(n1250) );
  and2 U1308 ( .A1(n539), .A2(n1247), .Z(n1249) );
  or2 U1309 ( .A1(n1250), .A2(n1249), .Z(n1251) );
  or2 U1310 ( .A1(n1252), .A2(n1251), .Z(n1253) );
  or2 U1312 ( .A1(n1255), .A2(n1256), .Z(n1264) );
  inv1 U1314 ( .I(n1256), .ZN(n1260) );
  or2 U1316 ( .A1(n1260), .A2(n1259), .Z(n1261) );
  or2 U1317 ( .A1(n1262), .A2(n1261), .Z(n1263) );
  or2 U1319 ( .A1(n1265), .A2(n1275), .Z(n1266) );
  and2 U1321 ( .A1(n1269), .A2(n1270), .Z(n1268) );
  inv1 U1322 ( .I(n1269), .ZN(n1271) );
  and2 U1323 ( .A1(n1271), .A2(n1270), .Z(n1273) );
  or2f U496 ( .A1(n1038), .A2(n757), .Z(n676) );
  inv1 U500 ( .I(n1054), .ZN(n1126) );
  or2f U501 ( .A1(n487), .A2(n1051), .Z(n1054) );
  and2 U502 ( .A1(h), .A2(n1007), .Z(n819) );
  inv1f U503 ( .I(j), .ZN(n1007) );
  inv1f U504 ( .I(n897), .ZN(n737) );
  and2 U505 ( .A1(n800), .A2(n799), .Z(n801) );
  or2 U506 ( .A1(n490), .A2(n1094), .Z(n754) );
  inv1 U507 ( .I(n773), .ZN(n868) );
  and2 U508 ( .A1(n816), .A2(n691), .Z(n475) );
  inv1 U509 ( .I(n1096), .ZN(n1097) );
  inv1 U510 ( .I(n523), .ZN(n668) );
  inv1 U512 ( .I(n1005), .ZN(n608) );
  and2 U513 ( .A1(n1233), .A2(n1232), .Z(n1244) );
  inv1 U515 ( .I(n752), .ZN(n1231) );
  inv1 U516 ( .I(n561), .ZN(n565) );
  or2 U518 ( .A1(n576), .A2(n543), .Z(n542) );
  or2 U519 ( .A1(n576), .A2(n580), .Z(n579) );
  inv1f U521 ( .I(n1058), .ZN(n540) );
  or2f U522 ( .A1(n955), .A2(y), .Z(n726) );
  or2f U524 ( .A1(n768), .A2(n591), .Z(n996) );
  inv1f U526 ( .I(n768), .ZN(n559) );
  inv1 U527 ( .I(n469), .ZN(n1196) );
  inv1f U529 ( .I(n664), .ZN(n518) );
  inv1f U532 ( .I(n), .ZN(n595) );
  or2f U537 ( .A1(n781), .A2(n634), .Z(n480) );
  inv1 U538 ( .I(n480), .ZN(n520) );
  or2f U539 ( .A1(n921), .A2(n922), .Z(n725) );
  or2f U542 ( .A1(n918), .A2(n922), .Z(n660) );
  inv1f U543 ( .I(n624), .ZN(n576) );
  inv1f U545 ( .I(n1233), .ZN(n769) );
  or2 U546 ( .A1(n656), .A2(n657), .Z(n790) );
  or2f U547 ( .A1(n782), .A2(n1234), .Z(n661) );
  or2f U548 ( .A1(n656), .A2(n1140), .Z(n633) );
  or2f U549 ( .A1(n710), .A2(n1234), .Z(n695) );
  inv1f U550 ( .I(n956), .ZN(n648) );
  inv1f U551 ( .I(n538), .ZN(n490) );
  and2f U553 ( .A1(n561), .A2(n1100), .Z(n1101) );
  or2f U555 ( .A1(n527), .A2(n839), .Z(n841) );
  inv1f U556 ( .I(n1085), .ZN(n1086) );
  and2f U558 ( .A1(n789), .A2(n1234), .Z(n657) );
  inv1f U560 ( .I(n766), .ZN(n789) );
  and2 U561 ( .A1(n857), .A2(b), .Z(n715) );
  inv1 U562 ( .I(n654), .ZN(n671) );
  or2 U563 ( .A1(n997), .A2(n883), .Z(n654) );
  and2 U564 ( .A1(n801), .A2(e), .Z(n802) );
  inv1 U565 ( .I(n707), .ZN(n793) );
  or2 U566 ( .A1(c), .A2(n975), .Z(n509) );
  and2 U567 ( .A1(n506), .A2(n858), .Z(n615) );
  inv1 U568 ( .I(n830), .ZN(n832) );
  inv1 U569 ( .I(w), .ZN(n875) );
  or2 U570 ( .A1(g0), .A2(n875), .Z(n885) );
  and2 U571 ( .A1(n1007), .A2(m), .Z(n892) );
  inv1 U573 ( .I(n727), .ZN(n915) );
  inv1 U574 ( .I(n508), .ZN(n815) );
  or2 U576 ( .A1(n700), .A2(n691), .Z(n628) );
  inv1 U577 ( .I(n476), .ZN(n973) );
  and2 U578 ( .A1(n524), .A2(n658), .Z(n656) );
  and2 U580 ( .A1(n577), .A2(n727), .Z(n584) );
  inv1 U582 ( .I(n582), .ZN(n771) );
  or2 U585 ( .A1(n915), .A2(n682), .Z(n483) );
  inv1 U586 ( .I(n907), .ZN(n909) );
  or2 U588 ( .A1(n1120), .A2(n511), .Z(n558) );
  and2 U589 ( .A1(n1093), .A2(n1117), .Z(n1118) );
  or2 U591 ( .A1(n1086), .A2(n622), .Z(n1117) );
  inv1 U592 ( .I(n743), .ZN(n989) );
  or2 U594 ( .A1(n757), .A2(n1057), .Z(n765) );
  inv1 U595 ( .I(n505), .ZN(n843) );
  or2 U596 ( .A1(n673), .A2(n672), .Z(n622) );
  inv1 U597 ( .I(n758), .ZN(n943) );
  or2 U598 ( .A1(n938), .A2(n940), .Z(n748) );
  and2 U599 ( .A1(n838), .A2(n837), .Z(n839) );
  or2 U601 ( .A1(n890), .A2(n889), .Z(n753) );
  or2 U602 ( .A1(n979), .A2(n553), .Z(n616) );
  or2 U604 ( .A1(n519), .A2(n518), .Z(n517) );
  or2 U606 ( .A1(n1036), .A2(n1023), .Z(n563) );
  or2 U608 ( .A1(n1039), .A2(n1080), .Z(n634) );
  or2 U610 ( .A1(n1221), .A2(n1220), .Z(n1225) );
  inv1 U611 ( .I(n725), .ZN(n923) );
  inv1 U615 ( .I(o), .ZN(n764) );
  inv1 U618 ( .I(g), .ZN(n1041) );
  inv1 U619 ( .I(h), .ZN(n528) );
  or2 U620 ( .A1(n1039), .A2(n1080), .Z(n1203) );
  or2 U621 ( .A1(n1080), .A2(n749), .Z(n1230) );
  inv1 U622 ( .I(n716), .ZN(n1153) );
  or2 U625 ( .A1(n1137), .A2(n1134), .Z(n1135) );
  or2 U629 ( .A1(n1172), .A2(n1171), .Z(a1) );
  inv1 U631 ( .I(n718), .ZN(n1172) );
  or2 U632 ( .A1(n1274), .A2(n610), .Z(f1) );
  or2 U634 ( .A1(n872), .A2(n687), .Z(n512) );
  or2 U636 ( .A1(n648), .A2(n1036), .Z(n651) );
  inv1f U638 ( .I(n535), .ZN(n659) );
  inv1 U639 ( .I(n969), .ZN(n1129) );
  or2f U641 ( .A1(n514), .A2(n932), .Z(n969) );
  inv1 U643 ( .I(n1047), .ZN(n1205) );
  inv1 U650 ( .I(n696), .ZN(n1020) );
  inv1 U652 ( .I(n692), .ZN(n696) );
  inv1 U653 ( .I(n513), .ZN(n646) );
  and2 U655 ( .A1(n528), .A2(e), .Z(n846) );
  or2 U656 ( .A1(n902), .A2(n903), .Z(n538) );
  or2f U661 ( .A1(n902), .A2(n903), .Z(n987) );
  and2 U663 ( .A1(n737), .A2(n889), .Z(n572) );
  and2f U664 ( .A1(n1014), .A2(j), .Z(n786) );
  and2f U665 ( .A1(n490), .A2(n1094), .Z(n561) );
  and2 U666 ( .A1(n1122), .A2(n768), .Z(n697) );
  or2f U667 ( .A1(n552), .A2(n768), .Z(n1024) );
  or2f U668 ( .A1(n864), .A2(n615), .Z(n867) );
  and2f U672 ( .A1(n1263), .A2(n1264), .Z(e1) );
  inv1 U675 ( .I(n1255), .ZN(n1262) );
  or2f U676 ( .A1(n741), .A2(n724), .Z(n488) );
  or2f U677 ( .A1(n973), .A2(n972), .Z(n544) );
  inv1 U678 ( .I(n920), .ZN(n922) );
  and2f U679 ( .A1(n909), .A2(n908), .Z(n910) );
  or2f U680 ( .A1(n473), .A2(n491), .Z(n787) );
  and2f U681 ( .A1(n916), .A2(n968), .Z(n618) );
  or2f U682 ( .A1(n475), .A2(n498), .Z(n481) );
  or2f U683 ( .A1(n592), .A2(n677), .Z(n524) );
  and2f U684 ( .A1(n863), .A2(n975), .Z(n756) );
  or2f U685 ( .A1(n637), .A2(n638), .Z(n1005) );
  or2f U686 ( .A1(n952), .A2(n668), .Z(n954) );
  or2f U687 ( .A1(n679), .A2(n1038), .Z(n1023) );
  and2 U689 ( .A1(n726), .A2(n953), .Z(n679) );
  or2f U693 ( .A1(n865), .A2(n777), .Z(n589) );
  or2f U695 ( .A1(n1128), .A2(n1127), .Z(n636) );
  or2f U698 ( .A1(n706), .A2(n568), .Z(n857) );
  or2f U700 ( .A1(n594), .A2(n1234), .Z(n706) );
  and2f U702 ( .A1(n735), .A2(n1234), .Z(n861) );
  and2f U704 ( .A1(n873), .A2(n1165), .Z(n743) );
  or2f U705 ( .A1(n1203), .A2(n1046), .Z(n1047) );
  or2f U706 ( .A1(n472), .A2(n601), .Z(n1046) );
  and2f U707 ( .A1(n880), .A2(n1234), .Z(n881) );
  or2f U708 ( .A1(n696), .A2(n1123), .Z(n1124) );
  or2f U709 ( .A1(n575), .A2(n490), .Z(n1019) );
  inv1f U710 ( .I(n591), .ZN(n575) );
  or2f U712 ( .A1(n494), .A2(n495), .Z(n813) );
  inv1f U714 ( .I(n704), .ZN(n814) );
  or2f U715 ( .A1(n548), .A2(n629), .Z(n627) );
  and2f U717 ( .A1(n886), .A2(n737), .Z(n573) );
  or2f U719 ( .A1(n501), .A2(n591), .Z(n1051) );
  and2f U720 ( .A1(n991), .A2(n990), .Z(n992) );
  inv1f U723 ( .I(n1006), .ZN(n607) );
  and2f U724 ( .A1(n509), .A2(n686), .Z(n807) );
  or2f U725 ( .A1(n604), .A2(n769), .Z(n603) );
  and2f U727 ( .A1(n635), .A2(n1140), .Z(n794) );
  or2f U728 ( .A1(n791), .A2(n790), .Z(n635) );
  or2f U731 ( .A1(n474), .A2(n690), .Z(n1233) );
  inv1f U732 ( .I(n529), .ZN(n673) );
  or2f U733 ( .A1(n530), .A2(n602), .Z(n529) );
  or2f U735 ( .A1(n885), .A2(n877), .Z(n831) );
  inv1f U736 ( .I(n553), .ZN(n530) );
  and2f U737 ( .A1(n554), .A2(n555), .Z(n599) );
  or2f U740 ( .A1(n955), .A2(y), .Z(n956) );
  inv1f U746 ( .I(n954), .ZN(n955) );
  and2f U747 ( .A1(n857), .A2(b), .Z(n506) );
  or2f U748 ( .A1(n1106), .A2(n1105), .Z(n1107) );
  or2f U750 ( .A1(n648), .A2(n676), .Z(n1096) );
  and2f U751 ( .A1(n1118), .A2(n697), .Z(n1223) );
  or2f U752 ( .A1(n1267), .A2(n1166), .Z(n1169) );
  or2f U754 ( .A1(n937), .A2(n748), .Z(n758) );
  or2f U755 ( .A1(n1004), .A2(n1019), .Z(n1006) );
  and2f U756 ( .A1(n716), .A2(n1150), .Z(n1156) );
  or2f U761 ( .A1(n803), .A2(n802), .Z(n907) );
  or2f U762 ( .A1(n1216), .A2(n1215), .Z(n1217) );
  or2f U764 ( .A1(n756), .A2(n583), .Z(n774) );
  and2f U766 ( .A1(n1231), .A2(n1247), .Z(n1232) );
  and2f U768 ( .A1(n956), .A2(n953), .Z(n522) );
  and2f U771 ( .A1(n1272), .A2(n1273), .Z(n1274) );
  or2f U772 ( .A1(n783), .A2(n1266), .Z(n1272) );
  or2f U773 ( .A1(n1269), .A2(n924), .Z(n925) );
  or2f U775 ( .A1(n705), .A2(n923), .Z(n1269) );
  or2f U776 ( .A1(n683), .A2(n681), .Z(n727) );
  or2f U777 ( .A1(n913), .A2(n1060), .Z(n683) );
  and2f U779 ( .A1(n858), .A2(n857), .Z(n859) );
  or2f U780 ( .A1(i), .A2(n855), .Z(n858) );
  and2f U782 ( .A1(n715), .A2(n858), .Z(n865) );
  or2f U788 ( .A1(n687), .A2(n751), .Z(n485) );
  or2f U789 ( .A1(n560), .A2(n1013), .Z(n477) );
  and2f U790 ( .A1(n537), .A2(n536), .Z(n903) );
  inv1f U791 ( .I(n736), .ZN(n536) );
  or2f U793 ( .A1(n754), .A2(n616), .Z(n1120) );
  and2f U798 ( .A1(n1178), .A2(n1179), .Z(n1180) );
  and2f U799 ( .A1(n873), .A2(n1165), .Z(n770) );
  inv1f U803 ( .I(n535), .ZN(n768) );
  and2f U806 ( .A1(n1170), .A2(n1169), .Z(n1171) );
  and2f U807 ( .A1(n713), .A2(n714), .Z(n810) );
  or2f U808 ( .A1(n803), .A2(n802), .Z(n713) );
  and2f U809 ( .A1(n933), .A2(n562), .Z(n714) );
  or2f U810 ( .A1(n688), .A2(n521), .Z(n933) );
  and2f U816 ( .A1(n1195), .A2(n1194), .Z(n1198) );
  and2f U817 ( .A1(n699), .A2(n700), .Z(n816) );
  or2f U818 ( .A1(n625), .A2(n712), .Z(n700) );
  and2f U820 ( .A1(n562), .A2(n933), .Z(n935) );
  or2f U821 ( .A1(n651), .A2(n676), .Z(n981) );
  or2f U823 ( .A1(n828), .A2(n827), .Z(n830) );
  and2f U824 ( .A1(n1032), .A2(c), .Z(n827) );
  or2f U825 ( .A1(n843), .A2(n842), .Z(n549) );
  and2f U826 ( .A1(n836), .A2(n835), .Z(n840) );
  or2f U827 ( .A1(n826), .A2(n825), .Z(n836) );
  and2f U828 ( .A1(n674), .A2(n873), .Z(n672) );
  and2f U829 ( .A1(n607), .A2(n608), .Z(n574) );
  or2f U830 ( .A1(n1169), .A2(n719), .Z(n718) );
  or2f U835 ( .A1(n649), .A2(n739), .Z(n1131) );
  or2f U836 ( .A1(n618), .A2(n617), .Z(n918) );
  and2f U837 ( .A1(n689), .A2(n619), .Z(n617) );
  or2f U839 ( .A1(n974), .A2(n981), .Z(n976) );
  or2f U841 ( .A1(n1018), .A2(n565), .Z(n974) );
  and2f U842 ( .A1(n584), .A2(n782), .Z(n916) );
  or2f U843 ( .A1(n508), .A2(e0), .Z(n625) );
  or2f U844 ( .A1(n794), .A2(n793), .Z(n508) );
  or2f U845 ( .A1(n646), .A2(g0), .Z(n1194) );
  and2f U847 ( .A1(n526), .A2(n1122), .Z(n1119) );
  and2f U848 ( .A1(n1093), .A2(n482), .Z(n526) );
  and2f U849 ( .A1(n879), .A2(i), .Z(n882) );
  inv1f U851 ( .I(n880), .ZN(n879) );
  or2f U854 ( .A1(n575), .A2(n518), .Z(n551) );
  and2f U856 ( .A1(n900), .A2(n901), .Z(n902) );
  or2f U865 ( .A1(n899), .A2(n670), .Z(n900) );
  and2f U866 ( .A1(n1187), .A2(n1188), .Z(n1189) );
  or2f U867 ( .A1(n783), .A2(n1183), .Z(n1187) );
  or2f U869 ( .A1(n680), .A2(n507), .Z(n873) );
  or2f U874 ( .A1(n871), .A2(e0), .Z(n680) );
  and2f U880 ( .A1(n863), .A2(n975), .Z(n864) );
  or2f U887 ( .A1(n862), .A2(n861), .Z(n863) );
  or2f U888 ( .A1(n1141), .A2(n691), .Z(n629) );
  or2f U889 ( .A1(n574), .A2(g0), .Z(n1221) );
  or2f U896 ( .A1(n471), .A2(n1018), .Z(n692) );
  or2f U898 ( .A1(n1128), .A2(n532), .Z(n1258) );
  and2f U899 ( .A1(n782), .A2(n935), .Z(n938) );
  or2f U902 ( .A1(n557), .A2(n1157), .Z(n953) );
  or2f U903 ( .A1(n468), .A2(n668), .Z(n557) );
  or2f U904 ( .A1(n929), .A2(z), .Z(n476) );
  or2f U910 ( .A1(n520), .A2(n1205), .Z(n484) );
  or2f U916 ( .A1(n911), .A2(n910), .Z(n920) );
  and2f U918 ( .A1(n759), .A2(n760), .Z(n1214) );
  inv1f U919 ( .I(n953), .ZN(n757) );
  or2 U920 ( .A1(n938), .A2(n937), .Z(n941) );
  or2f U921 ( .A1(n1053), .A2(n1087), .Z(n752) );
  or2f U923 ( .A1(n522), .A2(n1038), .Z(n1080) );
  inv1f U925 ( .I(n665), .ZN(n486) );
  or2f U926 ( .A1(n981), .A2(n982), .Z(n665) );
  or2f U930 ( .A1(n1267), .A2(n1174), .Z(n1178) );
  inv1f U932 ( .I(n775), .ZN(n1267) );
  and2f U934 ( .A1(n1154), .A2(n1153), .Z(n1155) );
  or2f U937 ( .A1(n1037), .A2(n1036), .Z(n1039) );
  inv1f U944 ( .I(n481), .ZN(n1037) );
  and2f U950 ( .A1(n775), .A2(n717), .Z(n716) );
  inv1f U954 ( .I(n712), .ZN(n1141) );
  or2f U958 ( .A1(n814), .A2(n813), .Z(n712) );
  or2f U959 ( .A1(n936), .A2(n669), .Z(n613) );
  or2f U960 ( .A1(n789), .A2(n788), .Z(n936) );
  and2f U961 ( .A1(n647), .A2(n934), .Z(n669) );
  and2f U963 ( .A1(n941), .A2(n940), .Z(n741) );
  or2f U964 ( .A1(n943), .A2(n488), .Z(n523) );
  and2f U965 ( .A1(n1247), .A2(n539), .Z(n545) );
  and2f U966 ( .A1(n540), .A2(n769), .Z(n539) );
  or2f U967 ( .A1(n648), .A2(n1038), .Z(n960) );
  or2f U970 ( .A1(n1178), .A2(n721), .Z(n720) );
  or2f U971 ( .A1(n1096), .A2(n994), .Z(n995) );
  or2f U972 ( .A1(n993), .A2(n992), .Z(n994) );
  or2f U973 ( .A1(n772), .A2(n771), .Z(n776) );
  and2f U979 ( .A1(n587), .A2(n588), .Z(n772) );
  inv1f U980 ( .I(n755), .ZN(n874) );
  or2f U981 ( .A1(n512), .A2(n751), .Z(n755) );
  inv1f U982 ( .I(n869), .ZN(n777) );
  or2f U983 ( .A1(n853), .A2(n852), .Z(n869) );
  or2f U990 ( .A1(n693), .A2(n1126), .Z(n532) );
  or2f U1000 ( .A1(n693), .A2(n1126), .Z(n1127) );
  or2f U1003 ( .A1(n1125), .A2(n1124), .Z(n1128) );
  or2f U1004 ( .A1(n1223), .A2(n1220), .Z(n1125) );
  or2f U1008 ( .A1(n478), .A2(n770), .Z(n1085) );
  or2f U1009 ( .A1(n553), .A2(n874), .Z(n478) );
  and2f U1012 ( .A1(n870), .A2(n777), .Z(n687) );
  or2f U1013 ( .A1(n868), .A2(n640), .Z(n870) );
  or2f U1014 ( .A1(n484), .A2(n497), .Z(n503) );
  or2f U1015 ( .A1(n484), .A2(n497), .Z(n534) );
  or2f U1017 ( .A1(n646), .A2(n486), .Z(n497) );
  or2f U1018 ( .A1(n673), .A2(n672), .Z(n778) );
  inv1f U1019 ( .I(n549), .ZN(n553) );
  or2f U1020 ( .A1(n549), .A2(a0), .Z(n504) );
  or2f U1023 ( .A1(n840), .A2(e0), .Z(n527) );
  and2f U1025 ( .A1(n830), .A2(n829), .Z(n834) );
  or2f U1026 ( .A1(n918), .A2(n919), .Z(n921) );
  inv1f U1027 ( .I(n550), .ZN(n919) );
  or2f U1028 ( .A1(n1207), .A2(n1131), .Z(n1133) );
  or2f U1029 ( .A1(n642), .A2(n1129), .Z(n1207) );
  or2f U1030 ( .A1(n917), .A2(n916), .Z(n1239) );
  and2f U1031 ( .A1(n689), .A2(n483), .Z(n917) );
  and2f U1043 ( .A1(n927), .A2(n928), .Z(n929) );
  and2f U1045 ( .A1(n926), .A2(n1275), .Z(n927) );
  and2f U1046 ( .A1(n921), .A2(n922), .Z(n705) );
  or2f U1047 ( .A1(n662), .A2(n878), .Z(n880) );
  and2f U1048 ( .A1(n663), .A2(n), .Z(n662) );
  and2f U1051 ( .A1(n711), .A2(p), .Z(n878) );
  or2f U1062 ( .A1(n1030), .A2(n563), .Z(n513) );
  or2f U1063 ( .A1(n603), .A2(n552), .Z(n1030) );
  or2f U1064 ( .A1(n1210), .A2(n1209), .Z(n626) );
  or2f U1068 ( .A1(n1202), .A2(n1201), .Z(n1210) );
  inv1f U1071 ( .I(n750), .ZN(n889) );
  or2f U1072 ( .A1(n671), .A2(n744), .Z(n750) );
  inv1f U1073 ( .I(n987), .ZN(n664) );
  or2f U1084 ( .A1(n575), .A2(n518), .Z(n552) );
  and2f U1085 ( .A1(n1258), .A2(n1257), .Z(n1259) );
  or2f U1089 ( .A1(n759), .A2(n1258), .Z(n1137) );
  or2f U1090 ( .A1(n1121), .A2(n559), .Z(n511) );
  or2f U1091 ( .A1(n765), .A2(n960), .Z(n493) );
  or2f U1092 ( .A1(n765), .A2(n960), .Z(n1121) );
  or2f U1102 ( .A1(n556), .A2(n937), .Z(n554) );
  or2f U1103 ( .A1(n938), .A2(e0), .Z(n556) );
  and2f U1109 ( .A1(n768), .A2(n1119), .Z(n763) );
  or2f U1115 ( .A1(n1254), .A2(n1253), .Z(n1255) );
  and2f U1118 ( .A1(n1229), .A2(n1228), .Z(n1254) );
  and2f U1121 ( .A1(n914), .A2(n1060), .Z(n682) );
  or2f U1127 ( .A1(n675), .A2(n912), .Z(n914) );
  and2f U1128 ( .A1(n930), .A2(n925), .Z(n591) );
  or2f U1132 ( .A1(n929), .A2(z), .Z(n930) );
  and2f U1133 ( .A1(n614), .A2(n1162), .Z(n1163) );
  or2f U1134 ( .A1(n576), .A2(n1158), .Z(n614) );
  or2f U1135 ( .A1(n1081), .A2(n490), .Z(n1040) );
  or2f U1141 ( .A1(n979), .A2(n553), .Z(n1081) );
  inv1f U1142 ( .I(n1011), .ZN(n979) );
  or2f U1143 ( .A1(n770), .A2(n874), .Z(n1011) );
  or2f U1147 ( .A1(n759), .A2(n1258), .Z(n624) );
  or2f U1149 ( .A1(n1133), .A2(n503), .Z(n759) );
  or2f U1150 ( .A1(n545), .A2(n606), .Z(n693) );
  and2f U1176 ( .A1(n607), .A2(n608), .Z(n606) );
  or2f U1182 ( .A1(n1211), .A2(n636), .Z(n775) );
  or2f U1183 ( .A1(n1133), .A2(n534), .Z(n1211) );
  or2f U1193 ( .A1(n474), .A2(n564), .Z(n535) );
  inv1f U1196 ( .I(n470), .ZN(n474) );
  or2f U1199 ( .A1(n789), .A2(n620), .Z(n782) );
  or2f U1205 ( .A1(n701), .A2(n1141), .Z(n699) );
endmodule

