
module C7552_iscas ( y6, x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, 
        k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, 
        s5, r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, 
        a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, 
        i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, 
        q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, 
        y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, h2, 
        g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, 
        o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, x0, 
        w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, 
        e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, 
        i, h, g, f, e, d, c, b, a, c11, b11, a11, z10, y10, x10, w10, v10, u10, 
        t10, s10, r10, q10, p10, o10, n10, m10, l10, k10, j10, i10, h10, g10, 
        f10, e10, d10, c10, b10, a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, 
        p9, o9, n9, m9, l9, k9, j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, 
        x8, w8, v8, u8, t8, s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, 
        f8, e8, d8, c8, b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, 
        n7, m7, l7, k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6 );
  input y6, x6, w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6,
         g6, f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, s5, r5, q5,
         p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5, z4,
         y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4,
         h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3,
         q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3,
         z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2,
         i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1,
         r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1,
         a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0,
         j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q,
         p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output c11, b11, a11, z10, y10, x10, w10, v10, u10, t10, s10, r10, q10, p10,
         o10, n10, m10, l10, k10, j10, i10, h10, g10, f10, e10, d10, c10, b10,
         a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9,
         j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8,
         s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8,
         b8, a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7,
         k7, j7, i7, h7, g7, f7, e7, d7, c7, b7, a7, z6;
  wire   w6, v6, u6, t6, s6, r6, q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6,
         f6, e6, d6, c6, b6, a6, z5, y5, x5, w5, v5, u5, t5, r5, q5, p5, o5,
         n5, m5, l5, i5, b1, a, x9, t9, y8, x8, n743, z850, n19, n118, n120,
         n121, n122, n124, n223, n224, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n403, n406, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n439, n456, n457,
         n458, n460, n463, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n529, n531, n535, n536, n537, n538, n553, n554, n555, n557, n560,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n628, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n643, n644,
         n657, n658, n659, n660, n661, n662, n663, n665, n666, n668, n669,
         n671, n672, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n711, n712, n713, n714, n715, n716, n717, n719, n720, n722, n723,
         n725, n726, n728, n729, n730, n731, n734, n737, n740, n741, n742,
         n744, n745, n746, n747, n748, n761, n762, n763, n764, n767, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n818, n819, n820, n821, n822, n824, n825, n826, n827,
         n828, n829, n832, n833, n834, n835, n836, n837, n838, n840, n841,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n868, n869, n870, n871, n872, n873, n874, n880,
         n885, n886, n887, n888, n889, n893, n895, n896, n897, n898, n900,
         n901, n902, n903, n904, n914, n915, n940, n941, n942, n943, n944,
         n945, n946, n947, n950, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n979, n990, n991, n996, n997, n998, n999, n1000,
         n1004, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1033, n1034, n1043, n1044, n1052, n1061, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1078, n1081, n1086,
         n1090, n1135, n1138, n1146, n1148, n1149, n1150, n1151, n1152, n1153,
         n1182, n1184, n1189, n1279, n1292, n1297, n1300, n1305, n1310, n1317,
         n1328, n1333, n1336, n1338, n1341, n1345, n1350, n1355, n1454, n1461,
         n1462, n1564, n1565, n1566, n1567, n1569, n1575, n1576, n1584, n1592,
         n1593, n1594, n1595, n1596, n1650, n1651, n1701, n1703, n1704, n1705,
         n1706, n1708, n1909, n1910, n1911, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1923, n1924, n1925, n1927, n1928, n1929,
         n1930, n1931, n1933, n1935, n1937, n1939, n1941, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2051, n2052, n2053, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2099, n2100, n2101, n2104,
         n2106, n2107, n2108, n2111, n2116, n2118, n2119, n2120, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         p10, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710;
  assign j8 = w6;
  assign i8 = v6;
  assign h8 = u6;
  assign g8 = t6;
  assign f8 = s6;
  assign e8 = r6;
  assign d8 = q6;
  assign c8 = p6;
  assign n8 = o6;
  assign b8 = n6;
  assign a8 = m6;
  assign z7 = l6;
  assign y7 = k6;
  assign x7 = j6;
  assign w7 = i6;
  assign v7 = h6;
  assign u7 = g6;
  assign t7 = f6;
  assign s7 = e6;
  assign r7 = d6;
  assign q7 = c6;
  assign p7 = b6;
  assign o7 = a6;
  assign n7 = z5;
  assign m7 = y5;
  assign l7 = x5;
  assign k7 = w5;
  assign j7 = v5;
  assign m8 = u5;
  assign i7 = t5;
  assign h7 = r5;
  assign g7 = q5;
  assign f7 = p5;
  assign e7 = o5;
  assign d7 = n5;
  assign l8 = m5;
  assign c7 = l5;
  assign z6 = i5;
  assign u8 = b1;
  assign a7 = a;
  assign b7 = a;
  assign t8 = a;
  assign b9 = a;
  assign h9 = x9;
  assign e9 = x9;
  assign h10 = x9;
  assign g9 = t9;
  assign f9 = t9;
  assign a9 = y8;
  assign v8 = x8;
  assign k8 = n743;
  assign w8 = n743;
  assign z8 = n743;
  assign n10 = z850;
  assign o10 = z850;
  assign q10 = p10;

  or2 U82 ( .A1(n120), .A2(n121), .Z(n118) );
  and2 U83 ( .A1(n122), .A2(n3659), .Z(n121) );
  and2 U84 ( .A1(n124), .A2(n3658), .Z(n120) );
  inv1 U161 ( .I(n223), .ZN(x8) );
  and2 U162 ( .A1(n224), .A2(j5), .Z(n223) );
  or2 U218 ( .A1(b), .A2(u), .Z(o8) );
  inv1 U227 ( .I(e), .ZN(n743) );
  or2 U304 ( .A1(n389), .A2(n390), .Z(g10) );
  or2 U305 ( .A1(p8), .A2(n391), .Z(n390) );
  or2 U306 ( .A1(q9), .A2(q8), .Z(n391) );
  inv1 U307 ( .I(n392), .ZN(q8) );
  and2 U308 ( .A1(n393), .A2(n394), .Z(n392) );
  and2 U309 ( .A1(l4), .A2(d4), .Z(n394) );
  and2 U310 ( .A1(x4), .A2(x1), .Z(n393) );
  or2 U311 ( .A1(n395), .A2(n396), .Z(q9) );
  or2 U312 ( .A1(n397), .A2(n398), .Z(n396) );
  or2 U313 ( .A1(n399), .A2(n400), .Z(n398) );
  inv1 U314 ( .I(n401), .ZN(n400) );
  or2 U315 ( .A1(n3660), .A2(n403), .Z(n401) );
  and2 U316 ( .A1(n403), .A2(n3660), .Z(n399) );
  and2 U323 ( .A1(n413), .A2(n414), .Z(n412) );
  or2 U324 ( .A1(n414), .A2(n413), .Z(n410) );
  or2 U325 ( .A1(n415), .A2(n416), .Z(n413) );
  and2 U326 ( .A1(n417), .A2(n418), .Z(n416) );
  inv1 U327 ( .I(n419), .ZN(n415) );
  or2 U328 ( .A1(n418), .A2(n417), .Z(n419) );
  or2 U353 ( .A1(n456), .A2(n457), .Z(n397) );
  inv1 U354 ( .I(n458), .ZN(n457) );
  or2 U355 ( .A1(n3661), .A2(n460), .Z(n458) );
  and2 U356 ( .A1(n460), .A2(n3661), .Z(n456) );
  and2 U361 ( .A1(n467), .A2(n468), .Z(n463) );
  and2 U363 ( .A1(n470), .A2(n471), .Z(n469) );
  or2 U364 ( .A1(n471), .A2(n470), .Z(n467) );
  or2 U365 ( .A1(n472), .A2(n473), .Z(n470) );
  and2 U366 ( .A1(n474), .A2(n475), .Z(n473) );
  inv1 U367 ( .I(n476), .ZN(n472) );
  or2 U368 ( .A1(n475), .A2(n474), .Z(n476) );
  or2 U394 ( .A1(n514), .A2(n515), .Z(n513) );
  and2 U395 ( .A1(n516), .A2(n517), .Z(n515) );
  inv1 U396 ( .I(n518), .ZN(n514) );
  or2 U397 ( .A1(n517), .A2(n516), .Z(n518) );
  or2 U398 ( .A1(n519), .A2(n520), .Z(n516) );
  and2 U407 ( .A1(f), .A2(n531), .Z(n529) );
  inv1 U408 ( .I(f4), .ZN(n531) );
  and2 U412 ( .A1(n535), .A2(n536), .Z(n517) );
  inv1 U413 ( .I(n537), .ZN(n536) );
  and2 U414 ( .A1(n538), .A2(n3662), .Z(n537) );
  or2 U415 ( .A1(n3662), .A2(n538), .Z(n535) );
  and2 U423 ( .A1(n553), .A2(n554), .Z(n512) );
  and2 U431 ( .A1(n564), .A2(n565), .Z(n560) );
  and2 U433 ( .A1(n567), .A2(n568), .Z(n566) );
  or2 U434 ( .A1(n568), .A2(n567), .Z(n564) );
  or2 U435 ( .A1(n569), .A2(n570), .Z(n567) );
  and2 U436 ( .A1(n571), .A2(n572), .Z(n570) );
  inv1 U437 ( .I(n573), .ZN(n569) );
  or2 U438 ( .A1(n572), .A2(n571), .Z(n573) );
  or2 U439 ( .A1(n574), .A2(n575), .Z(n571) );
  inv1 U463 ( .I(n608), .ZN(p8) );
  and2 U464 ( .A1(n609), .A2(n610), .Z(n608) );
  and2 U465 ( .A1(h5), .A2(d3), .Z(n610) );
  and2 U466 ( .A1(v4), .A2(v1), .Z(n609) );
  or2 U467 ( .A1(n611), .A2(n612), .Z(n389) );
  inv1 U469 ( .I(n613), .ZN(r8) );
  and2 U470 ( .A1(n614), .A2(n615), .Z(n613) );
  and2 U471 ( .A1(c3), .A2(b3), .Z(n615) );
  and2 U472 ( .A1(f3), .A2(e3), .Z(n614) );
  or2 U475 ( .A1(n620), .A2(n621), .Z(n619) );
  inv1 U476 ( .I(n622), .ZN(n621) );
  and2 U478 ( .A1(n624), .A2(n623), .Z(n620) );
  or2 U485 ( .A1(n633), .A2(n634), .Z(n632) );
  and2 U486 ( .A1(n634), .A2(n633), .Z(n630) );
  and2 U489 ( .A1(n638), .A2(n639), .Z(n637) );
  or2 U490 ( .A1(n639), .A2(n638), .Z(n635) );
  or2 U491 ( .A1(n640), .A2(n641), .Z(n638) );
  and2 U492 ( .A1(n3664), .A2(n643), .Z(n641) );
  and2 U494 ( .A1(n3665), .A2(n644), .Z(n640) );
  or2 U507 ( .A1(n657), .A2(n658), .Z(n634) );
  and2 U508 ( .A1(n659), .A2(n660), .Z(n658) );
  inv1 U509 ( .I(n661), .ZN(n657) );
  or2 U510 ( .A1(n659), .A2(n660), .Z(n661) );
  or2 U511 ( .A1(n662), .A2(n663), .Z(n659) );
  and2 U512 ( .A1(n3666), .A2(n665), .Z(n663) );
  and2 U514 ( .A1(n3667), .A2(n666), .Z(n662) );
  or2 U516 ( .A1(n668), .A2(n669), .Z(n624) );
  and2 U517 ( .A1(n3668), .A2(n671), .Z(n669) );
  and2 U519 ( .A1(n3669), .A2(n672), .Z(n668) );
  or2 U521 ( .A1(n674), .A2(n675), .Z(n618) );
  inv1 U522 ( .I(n676), .ZN(n675) );
  and2 U524 ( .A1(n678), .A2(n677), .Z(n674) );
  or2 U528 ( .A1(n682), .A2(n683), .Z(n679) );
  and2 U530 ( .A1(n686), .A2(n687), .Z(n685) );
  inv1 U531 ( .I(n688), .ZN(n684) );
  or2 U532 ( .A1(n687), .A2(n686), .Z(n688) );
  or2 U533 ( .A1(n689), .A2(n690), .Z(n686) );
  and2 U534 ( .A1(n691), .A2(n692), .Z(n690) );
  inv1 U535 ( .I(n693), .ZN(n689) );
  or2 U536 ( .A1(n692), .A2(n691), .Z(n693) );
  and2 U553 ( .A1(n711), .A2(n712), .Z(n687) );
  inv1 U554 ( .I(n713), .ZN(n712) );
  and2 U555 ( .A1(n714), .A2(n715), .Z(n713) );
  or2 U556 ( .A1(n714), .A2(n715), .Z(n711) );
  or2 U557 ( .A1(n716), .A2(n717), .Z(n714) );
  and2 U558 ( .A1(n3670), .A2(n719), .Z(n717) );
  inv1 U559 ( .I(n720), .ZN(n716) );
  or2 U560 ( .A1(n719), .A2(n3670), .Z(n720) );
  or2 U562 ( .A1(n722), .A2(n723), .Z(n678) );
  and2 U563 ( .A1(n3671), .A2(n725), .Z(n723) );
  and2 U565 ( .A1(n3672), .A2(n726), .Z(n722) );
  and2 U569 ( .A1(n3673), .A2(n3674), .Z(n731) );
  inv1 U570 ( .I(n734), .ZN(n730) );
  and2 U577 ( .A1(n742), .A2(n744), .Z(n741) );
  inv1 U581 ( .I(n748), .ZN(n747) );
  or2 U582 ( .A1(n3675), .A2(n3676), .Z(n748) );
  and2 U583 ( .A1(n3676), .A2(n3675), .Z(n746) );
  and2 U592 ( .A1(f), .A2(n762), .Z(n761) );
  or2 U593 ( .A1(n763), .A2(n764), .Z(n762) );
  and2 U594 ( .A1(n3677), .A2(n2580), .Z(n764) );
  and2 U596 ( .A1(e6), .A2(n767), .Z(n763) );
  and2 U619 ( .A1(n790), .A2(n791), .Z(n728) );
  or2 U620 ( .A1(n792), .A2(n793), .Z(n791) );
  inv1 U621 ( .I(n794), .ZN(n790) );
  and2 U622 ( .A1(n793), .A2(n792), .Z(n794) );
  or2 U623 ( .A1(n795), .A2(n796), .Z(n792) );
  and2 U624 ( .A1(n797), .A2(n798), .Z(n796) );
  inv1 U625 ( .I(n799), .ZN(n795) );
  or2 U626 ( .A1(n798), .A2(n797), .Z(n799) );
  or2 U627 ( .A1(n800), .A2(n801), .Z(n797) );
  and2 U628 ( .A1(n802), .A2(n803), .Z(n801) );
  and2 U630 ( .A1(n3681), .A2(n804), .Z(n800) );
  and2 U632 ( .A1(f), .A2(n808), .Z(n807) );
  or2 U633 ( .A1(n809), .A2(n810), .Z(n808) );
  inv1 U634 ( .I(n811), .ZN(n810) );
  or2 U635 ( .A1(n812), .A2(l5), .Z(n811) );
  and2 U636 ( .A1(l5), .A2(n812), .Z(n809) );
  and2 U638 ( .A1(n814), .A2(n815), .Z(n813) );
  and2 U640 ( .A1(n812), .A2(h1), .Z(n816) );
  or2 U641 ( .A1(h1), .A2(n812), .Z(n814) );
  and2 U644 ( .A1(f), .A2(n819), .Z(n818) );
  or2 U645 ( .A1(n820), .A2(n821), .Z(n819) );
  inv1 U646 ( .I(n822), .ZN(n821) );
  or2 U647 ( .A1(n3701), .A2(r5), .Z(n822) );
  and2 U648 ( .A1(r5), .A2(n3701), .Z(n820) );
  and2 U650 ( .A1(n825), .A2(n826), .Z(n824) );
  or2 U651 ( .A1(n827), .A2(n828), .Z(n826) );
  or2 U652 ( .A1(s5), .A2(n3701), .Z(n825) );
  or2 U656 ( .A1(n3698), .A2(f), .Z(n829) );
  and2 U657 ( .A1(n832), .A2(n833), .Z(n793) );
  inv1 U658 ( .I(n834), .ZN(n833) );
  and2 U659 ( .A1(n835), .A2(n836), .Z(n834) );
  or2 U660 ( .A1(n835), .A2(n836), .Z(n832) );
  or2 U661 ( .A1(n837), .A2(n838), .Z(n835) );
  and2 U662 ( .A1(n3680), .A2(n840), .Z(n838) );
  and2 U664 ( .A1(n3678), .A2(n841), .Z(n837) );
  or2 U666 ( .A1(s9), .A2(s8), .Z(n611) );
  inv1 U667 ( .I(n843), .ZN(s8) );
  and2 U668 ( .A1(n844), .A2(n845), .Z(n843) );
  and2 U669 ( .A1(h3), .A2(h2), .Z(n845) );
  and2 U670 ( .A1(s3), .A2(r2), .Z(n844) );
  or2 U673 ( .A1(n850), .A2(n851), .Z(n849) );
  and2 U674 ( .A1(n852), .A2(n853), .Z(n851) );
  inv1 U675 ( .I(n854), .ZN(n850) );
  or2 U676 ( .A1(n853), .A2(n852), .Z(n854) );
  or2 U677 ( .A1(n855), .A2(n856), .Z(n852) );
  and2 U691 ( .A1(n868), .A2(n869), .Z(n853) );
  inv1 U692 ( .I(n870), .ZN(n869) );
  and2 U693 ( .A1(n871), .A2(n872), .Z(n870) );
  or2 U694 ( .A1(n872), .A2(n871), .Z(n868) );
  or2 U695 ( .A1(n873), .A2(n874), .Z(n871) );
  and2 U700 ( .A1(n3702), .A2(n880), .Z(n872) );
  or2 U705 ( .A1(n885), .A2(n886), .Z(n848) );
  inv1 U706 ( .I(n887), .ZN(n886) );
  and2 U708 ( .A1(n889), .A2(n888), .Z(n885) );
  or2 U720 ( .A1(n904), .A2(n903), .Z(n900) );
  and2 U728 ( .A1(n915), .A2(f), .Z(n914) );
  inv1 U737 ( .I(n), .ZN(n439) );
  or2 U753 ( .A1(n942), .A2(n943), .Z(n941) );
  inv1 U754 ( .I(n944), .ZN(n943) );
  or2 U761 ( .A1(n952), .A2(n953), .Z(n950) );
  and2 U762 ( .A1(n954), .A2(n955), .Z(n953) );
  inv1 U763 ( .I(n956), .ZN(n952) );
  or2 U764 ( .A1(n955), .A2(n954), .Z(n956) );
  or2 U765 ( .A1(n957), .A2(n958), .Z(n954) );
  and2 U766 ( .A1(n959), .A2(n960), .Z(n958) );
  inv1 U767 ( .I(n961), .ZN(n957) );
  or2 U768 ( .A1(n960), .A2(n959), .Z(n961) );
  and2 U785 ( .A1(n979), .A2(n3704), .Z(n955) );
  or2 U794 ( .A1(n990), .A2(n991), .Z(n946) );
  inv1 U800 ( .I(n998), .ZN(n997) );
  or2 U802 ( .A1(n1000), .A2(n999), .Z(n996) );
  inv1 U808 ( .I(n1008), .ZN(n1007) );
  inv1 U812 ( .I(n1013), .ZN(n1012) );
  and2 U813 ( .A1(n1014), .A2(n1015), .Z(n1013) );
  or2 U814 ( .A1(n1015), .A2(n1014), .Z(n1011) );
  or2 U815 ( .A1(n1016), .A2(n1017), .Z(n1014) );
  or2 U831 ( .A1(n1033), .A2(n1034), .Z(n1010) );
  or2 U839 ( .A1(n1043), .A2(n1044), .Z(n1000) );
  and2 U854 ( .A1(n1063), .A2(n1064), .Z(n1061) );
  or2 U855 ( .A1(n1065), .A2(n1066), .Z(n1064) );
  and2 U857 ( .A1(n1067), .A2(n1068), .Z(n1065) );
  or2 U858 ( .A1(n1069), .A2(n1070), .Z(n1068) );
  and2 U867 ( .A1(f), .A2(n3696), .Z(n1078) );
  and2 U874 ( .A1(f), .A2(n3699), .Z(n1081) );
  and2 U880 ( .A1(f), .A2(n3695), .Z(n1086) );
  and2 U886 ( .A1(f), .A2(n3694), .Z(n1090) );
  and2 U921 ( .A1(f), .A2(n3692), .Z(n1135) );
  and2 U924 ( .A1(x2), .A2(f), .Z(n1138) );
  and2 U932 ( .A1(n1148), .A2(n1149), .Z(n1146) );
  or2 U933 ( .A1(n1150), .A2(n1151), .Z(n1149) );
  and2 U935 ( .A1(n1152), .A2(n1153), .Z(n1150) );
  and2 U960 ( .A1(m3), .A2(f), .Z(n1182) );
  and2 U963 ( .A1(n3), .A2(f), .Z(n1184) );
  and2 U970 ( .A1(o3), .A2(f), .Z(n1189) );
  and2 U1064 ( .A1(t3), .A2(f), .Z(n1279) );
  and2 U1078 ( .A1(l3), .A2(f), .Z(n1292) );
  and2 U1084 ( .A1(f), .A2(n3686), .Z(n1297) );
  and2 U1087 ( .A1(i3), .A2(f), .Z(n1300) );
  and2 U1094 ( .A1(j3), .A2(f), .Z(n1305) );
  and2 U1100 ( .A1(k3), .A2(f), .Z(n1310) );
  and2 U1110 ( .A1(f), .A2(n3691), .Z(n1317) );
  and2 U1125 ( .A1(f), .A2(n3688), .Z(n1328) );
  and2 U1134 ( .A1(y2), .A2(n2107), .Z(n1336) );
  and2 U1137 ( .A1(f), .A2(n3690), .Z(n1338) );
  and2 U1146 ( .A1(f), .A2(n3689), .Z(n1341) );
  and2 U1152 ( .A1(f), .A2(n3687), .Z(n1345) );
  and2 U1157 ( .A1(f), .A2(n3697), .Z(n1350) );
  and2 U1162 ( .A1(n3698), .A2(n3700), .Z(n1355) );
  and2 U1165 ( .A1(n828), .A2(y6), .Z(n1052) );
  inv1 U1166 ( .I(s5), .ZN(n828) );
  and2 U1190 ( .A1(i2), .A2(a), .Z(c9) );
  or2 U1265 ( .A1(n1461), .A2(n1462), .Z(n1454) );
  or2 U1362 ( .A1(n1565), .A2(n1566), .Z(n1564) );
  or2 U1364 ( .A1(n3682), .A2(n1569), .Z(n1567) );
  and2 U1365 ( .A1(n1569), .A2(n3682), .Z(n1565) );
  or2 U1371 ( .A1(n1575), .A2(n1576), .Z(n1569) );
  or2 U1394 ( .A1(n1592), .A2(n1593), .Z(n1584) );
  and2 U1395 ( .A1(n1594), .A2(n1595), .Z(n1593) );
  and2 U1397 ( .A1(n1596), .A2(n3683), .Z(n1592) );
  inv1 U1462 ( .I(n1650), .ZN(y8) );
  and2 U1463 ( .A1(n1651), .A2(p1), .Z(n1650) );
  and2 U1464 ( .A1(o1), .A2(n224), .Z(n1651) );
  inv1 U1465 ( .I(b), .ZN(n224) );
  or2 U1512 ( .A1(n1703), .A2(n1704), .Z(n1701) );
  and2 U1513 ( .A1(n19), .A2(n3705), .Z(n1704) );
  and2 U1515 ( .A1(n3685), .A2(n3684), .Z(n1703) );
  and2 U1518 ( .A1(n1706), .A2(n3700), .Z(n1705) );
  and2 U1521 ( .A1(y6), .A2(r5), .Z(n1706) );
  and2 U1528 ( .A1(q5), .A2(y6), .Z(n1708) );
  or2 U1955 ( .A1(n2496), .A2(n1925), .Z(n1909) );
  inv1 U1958 ( .I(n2065), .ZN(n1911) );
  and2 U1960 ( .A1(n1970), .A2(n2290), .Z(n1913) );
  and2 U1961 ( .A1(n3209), .A2(n3212), .Z(n1914) );
  inv1 U1962 ( .I(n1914), .ZN(n3214) );
  inv1 U1966 ( .I(n3051), .ZN(n1918) );
  inv1 U1969 ( .I(n1920), .ZN(n2058) );
  and2 U1970 ( .A1(n1946), .A2(u1), .Z(n1921) );
  and2 U1973 ( .A1(n1946), .A2(n1), .Z(n1924) );
  and2 U1974 ( .A1(n2049), .A2(j1), .Z(n1925) );
  and2 U1976 ( .A1(n1946), .A2(a1), .Z(n1927) );
  and2 U1978 ( .A1(n3710), .A2(g), .Z(n1929) );
  and2 U1982 ( .A1(n2119), .A2(d0), .Z(n1933) );
  and2 U1984 ( .A1(n2111), .A2(k1), .Z(n1935) );
  and2 U1986 ( .A1(n2111), .A2(x0), .Z(n1937) );
  and2 U1988 ( .A1(n2122), .A2(z0), .Z(n1939) );
  and2 U1990 ( .A1(n2116), .A2(t1), .Z(n1941) );
  and2 U1992 ( .A1(n2049), .A2(q1), .Z(n1943) );
  and2 U1996 ( .A1(n1946), .A2(k), .Z(n1947) );
  and2 U1997 ( .A1(n1946), .A2(y0), .Z(n1948) );
  and2 U2002 ( .A1(n2025), .A2(n2084), .Z(n1953) );
  inv1 U2003 ( .I(n1953), .ZN(n2026) );
  inv1 U2005 ( .I(n2078), .ZN(n1955) );
  and2 U2008 ( .A1(n2032), .A2(n2033), .Z(n1957) );
  and2 U2009 ( .A1(n2905), .A2(n2032), .Z(n1958) );
  and2 U2011 ( .A1(n1959), .A2(n1960), .Z(n2827) );
  or2 U2012 ( .A1(n2826), .A2(n2030), .Z(n1960) );
  or2 U2013 ( .A1(n2031), .A2(n2826), .Z(n1961) );
  inv1 U2015 ( .I(n1962), .ZN(n2125) );
  or2 U2017 ( .A1(n2458), .A2(n2636), .Z(n1964) );
  and2 U2018 ( .A1(n1966), .A2(n2221), .Z(n1965) );
  inv1 U2019 ( .I(n1965), .ZN(n2637) );
  inv1 U2020 ( .I(n2458), .ZN(n1966) );
  or2 U2021 ( .A1(n1968), .A2(n3612), .Z(n1967) );
  and2 U2023 ( .A1(n1970), .A2(n2290), .Z(n1969) );
  inv1 U2025 ( .I(n2569), .ZN(n1970) );
  or2 U2026 ( .A1(n3062), .A2(n1971), .Z(n2040) );
  and2 U2028 ( .A1(n3005), .A2(n2019), .Z(n1972) );
  and2 U2029 ( .A1(n2085), .A2(n2160), .Z(n1973) );
  inv1 U2030 ( .I(n1973), .ZN(n1974) );
  or2 U2032 ( .A1(n2943), .A2(n2027), .Z(n1975) );
  or2 U2033 ( .A1(n3061), .A2(n1978), .Z(n1976) );
  or2 U2035 ( .A1(n3446), .A2(n1955), .Z(n1977) );
  or2 U2036 ( .A1(n3062), .A2(n3446), .Z(n1978) );
  inv1 U2041 ( .I(n2670), .ZN(n1982) );
  inv1 U2043 ( .I(n1983), .ZN(n3152) );
  and2 U2044 ( .A1(n2626), .A2(n2625), .Z(n1984) );
  and2 U2045 ( .A1(n2045), .A2(n2125), .Z(n1985) );
  or2 U2053 ( .A1(n3360), .A2(n3359), .Z(n1991) );
  and2 U2055 ( .A1(n3370), .A2(n3358), .Z(n1993) );
  or2 U2056 ( .A1(n1993), .A2(n1994), .Z(n3365) );
  and2 U2058 ( .A1(n1996), .A2(n2603), .Z(n1995) );
  inv1 U2059 ( .I(n1995), .ZN(n3458) );
  inv1 U2060 ( .I(n2604), .ZN(n1996) );
  inv1 U2061 ( .I(n3370), .ZN(n1997) );
  and2 U2062 ( .A1(n3630), .A2(n3629), .Z(n1999) );
  and2 U2068 ( .A1(n3508), .A2(n2006), .Z(n2004) );
  or2 U2073 ( .A1(n3484), .A2(n2008), .Z(n2007) );
  inv1 U2074 ( .I(n3466), .ZN(n2008) );
  or2 U2075 ( .A1(n2138), .A2(n3139), .Z(n2009) );
  or2 U2076 ( .A1(n1984), .A2(n3242), .Z(n2010) );
  or2 U2077 ( .A1(n2649), .A2(n2013), .Z(n2011) );
  or2 U2079 ( .A1(n2092), .A2(n2093), .Z(n2012) );
  or2 U2080 ( .A1(n2648), .A2(n2092), .Z(n2013) );
  or2 U2082 ( .A1(n2434), .A2(n1921), .Z(n2015) );
  and2 U2083 ( .A1(n2672), .A2(n1955), .Z(n2016) );
  inv1 U2085 ( .I(g6), .ZN(n2018) );
  inv1 U2087 ( .I(n2019), .ZN(n3201) );
  inv1 U2088 ( .I(n2632), .ZN(n2020) );
  inv1 U2090 ( .I(n2021), .ZN(n3441) );
  and2 U2095 ( .A1(n2085), .A2(n2160), .Z(n2025) );
  inv1 U2096 ( .I(n2084), .ZN(n2027) );
  and2 U2097 ( .A1(n2153), .A2(n2100), .Z(n2028) );
  or2 U2100 ( .A1(n2825), .A2(n2824), .Z(n2030) );
  or2 U2101 ( .A1(n2822), .A2(n2825), .Z(n2031) );
  or2 U2102 ( .A1(n2916), .A2(n2915), .Z(n2032) );
  or2 U2103 ( .A1(n2914), .A2(n2916), .Z(n2033) );
  inv1 U2106 ( .I(n2034), .ZN(n3119) );
  and2 U2107 ( .A1(n1995), .A2(n2008), .Z(n2036) );
  and2 U2108 ( .A1(n1988), .A2(n1995), .Z(n2037) );
  or2 U2109 ( .A1(n2034), .A2(n3491), .Z(n2038) );
  inv1 U2110 ( .I(n2038), .ZN(n2066) );
  inv1 U2112 ( .I(n2040), .ZN(n2039) );
  or2 U2115 ( .A1(n2126), .A2(n2172), .Z(n2043) );
  and2 U2116 ( .A1(n2045), .A2(n2125), .Z(n2044) );
  inv1 U2117 ( .I(n1985), .ZN(n2514) );
  inv1 U2118 ( .I(n2126), .ZN(n2045) );
  or2 U2119 ( .A1(n2048), .A2(n2046), .Z(n2991) );
  inv1 U2122 ( .I(n2047), .ZN(n2064) );
  and2 U2127 ( .A1(n2051), .A2(n2052), .Z(n3050) );
  or2 U2128 ( .A1(n3355), .A2(n2595), .Z(n2052) );
  or2 U2129 ( .A1(n3313), .A2(n3355), .Z(n2053) );
  inv1 U2133 ( .I(n2056), .ZN(n2057) );
  inv1 U2138 ( .I(n2062), .ZN(n3095) );
  and2 U2139 ( .A1(n3309), .A2(n2695), .Z(n2063) );
  and2 U2141 ( .A1(n2634), .A2(n2633), .Z(n2067) );
  inv1 U2142 ( .I(n2014), .ZN(n3230) );
  inv1 U2144 ( .I(n2068), .ZN(n3191) );
  inv1 U2145 ( .I(n2642), .ZN(n2069) );
  and2 U2146 ( .A1(n2088), .A2(n2658), .Z(n2070) );
  or2 U2149 ( .A1(n2161), .A2(n2073), .Z(n2086) );
  inv1 U2151 ( .I(n3467), .ZN(n2074) );
  and2 U2152 ( .A1(n3494), .A2(n2077), .Z(n2075) );
  and2 U2154 ( .A1(n1995), .A2(n2614), .Z(n2076) );
  and2 U2163 ( .A1(n2595), .A2(n3355), .Z(n2083) );
  and2 U2165 ( .A1(n2084), .A2(n2085), .Z(n2163) );
  and2 U2167 ( .A1(n2088), .A2(n2658), .Z(n2087) );
  inv1 U2169 ( .I(n2659), .ZN(n2088) );
  and2 U2170 ( .A1(n2090), .A2(n2256), .Z(n2089) );
  inv1 U2171 ( .I(n2089), .ZN(n2581) );
  inv1 U2172 ( .I(n2536), .ZN(n2090) );
  inv1 U2173 ( .I(n1915), .ZN(n2957) );
  or2 U2174 ( .A1(n2667), .A2(n2017), .Z(n2091) );
  and2 U2177 ( .A1(n2019), .A2(n3189), .Z(n2093) );
  inv1 U2179 ( .I(n1972), .ZN(n3007) );
  and2 U2182 ( .A1(n2960), .A2(n2157), .Z(n2097) );
  inv1 U2183 ( .I(n2097), .ZN(n2162) );
  and2 U2185 ( .A1(n2153), .A2(n2100), .Z(n2099) );
  inv1 U2186 ( .I(n2028), .ZN(n3531) );
  inv1 U2187 ( .I(n2154), .ZN(n2100) );
  inv1 U2203 ( .I(f), .ZN(n2116) );
  inv1 U2210 ( .I(l), .ZN(n3700) );
  or2 U2211 ( .A1(n3700), .A2(n1708), .Z(n3705) );
  inv1 U2212 ( .I(n3705), .ZN(n3685) );
  or2 U2213 ( .A1(n3700), .A2(n1706), .Z(n2123) );
  inv1 U2214 ( .I(n2123), .ZN(n2716) );
  or2 U2215 ( .A1(n2716), .A2(n1705), .Z(n19) );
  inv1 U2216 ( .I(n19), .ZN(n3684) );
  and2 U2217 ( .A1(p4), .A2(f), .Z(n2124) );
  inv1 U2219 ( .I(n2507), .ZN(n2509) );
  and2 U2220 ( .A1(o4), .A2(f), .Z(n2126) );
  inv1 U2221 ( .I(u6), .ZN(n2172) );
  or2 U2222 ( .A1(n2043), .A2(n1962), .Z(n2140) );
  inv1 U2227 ( .I(n2143), .ZN(n3145) );
  and2 U2228 ( .A1(n3152), .A2(n3145), .Z(n2130) );
  and2 U2229 ( .A1(n1983), .A2(n2143), .Z(n2129) );
  or2 U2230 ( .A1(n2130), .A2(n2129), .Z(n1596) );
  and2 U2231 ( .A1(n4), .A2(n2106), .Z(n2131) );
  or2 U2232 ( .A1(n2131), .A2(n1952), .Z(n2512) );
  inv1 U2233 ( .I(n2512), .ZN(n2513) );
  and2 U2234 ( .A1(v6), .A2(n2513), .Z(n2133) );
  or2 U2235 ( .A1(n2513), .A2(v6), .Z(n2132) );
  and2 U2241 ( .A1(m4), .A2(f), .Z(n2135) );
  or2 U2242 ( .A1(n2135), .A2(n1933), .Z(n2518) );
  inv1 U2243 ( .I(n2518), .ZN(n2520) );
  and2 U2244 ( .A1(w6), .A2(n2520), .Z(n2136) );
  or2 U2245 ( .A1(n2520), .A2(w6), .Z(n2625) );
  inv1 U2246 ( .I(n2625), .ZN(n2696) );
  inv1 U2248 ( .I(n3139), .ZN(n3136) );
  or2 U2249 ( .A1(n2137), .A2(n3136), .Z(n2147) );
  inv1 U2250 ( .I(n2147), .ZN(n2139) );
  inv1 U2251 ( .I(n2137), .ZN(n2138) );
  inv1 U2253 ( .I(n2009), .ZN(n2697) );
  or2 U2254 ( .A1(n2139), .A2(n2697), .Z(n1594) );
  inv1 U2255 ( .I(n1594), .ZN(n3683) );
  inv1 U2256 ( .I(n1596), .ZN(n1595) );
  inv1 U2257 ( .I(t6), .ZN(n2169) );
  or2 U2258 ( .A1(n2507), .A2(n2169), .Z(n3156) );
  inv1 U2259 ( .I(n3156), .ZN(n3158) );
  inv1 U2260 ( .I(n2140), .ZN(n2142) );
  or2 U2261 ( .A1(n2142), .A2(n2141), .Z(n3426) );
  inv1 U2262 ( .I(n3426), .ZN(n3423) );
  or2 U2263 ( .A1(n3158), .A2(n1983), .Z(n3417) );
  inv1 U2264 ( .I(n3417), .ZN(n3419) );
  and2 U2265 ( .A1(n3423), .A2(n3419), .Z(n2144) );
  or2 U2266 ( .A1(n2144), .A2(n2143), .Z(n3133) );
  and2 U2267 ( .A1(n3158), .A2(n3133), .Z(n1575) );
  inv1 U2268 ( .I(n3133), .ZN(n3146) );
  and2 U2269 ( .A1(n3156), .A2(n3146), .Z(n1576) );
  inv1 U2272 ( .I(n2623), .ZN(n2146) );
  and2 U2273 ( .A1(n3139), .A2(n2146), .Z(n2149) );
  and2 U2274 ( .A1(n2147), .A2(n2623), .Z(n2148) );
  or2 U2275 ( .A1(n2149), .A2(n2148), .Z(n2150) );
  and2 U2276 ( .A1(n2150), .A2(n2009), .Z(n3682) );
  inv1 U2277 ( .I(n1567), .ZN(n1566) );
  and2 U2278 ( .A1(b5), .A2(n2079), .Z(n2151) );
  or2 U2279 ( .A1(n2058), .A2(j6), .Z(n2970) );
  and2 U2281 ( .A1(a5), .A2(f), .Z(n2152) );
  or2 U2284 ( .A1(n2549), .A2(k6), .Z(n2153) );
  and2 U2285 ( .A1(k6), .A2(n2549), .Z(n2154) );
  and2 U2286 ( .A1(n2969), .A2(n2099), .Z(n2155) );
  and2 U2287 ( .A1(z4), .A2(n2106), .Z(n2156) );
  and2 U2290 ( .A1(l6), .A2(n2559), .Z(n2158) );
  and2 U2294 ( .A1(y4), .A2(f), .Z(n2159) );
  or2 U2295 ( .A1(n2159), .A2(n1939), .Z(n2553) );
  inv1 U2296 ( .I(n2553), .ZN(n2552) );
  and2 U2297 ( .A1(m6), .A2(n2552), .Z(n2161) );
  or2 U2298 ( .A1(n2552), .A2(m6), .Z(n2160) );
  inv1 U2299 ( .I(n2160), .ZN(n2619) );
  inv1 U2301 ( .I(n3554), .ZN(n2949) );
  or2 U2302 ( .A1(n2162), .A2(n2949), .Z(n3551) );
  inv1 U2303 ( .I(n2163), .ZN(n3559) );
  or2 U2304 ( .A1(n3552), .A2(n3559), .Z(n2168) );
  inv1 U2305 ( .I(n2168), .ZN(n2944) );
  and2 U2306 ( .A1(n2970), .A2(n1915), .Z(n2165) );
  and2 U2307 ( .A1(n2969), .A2(n2957), .Z(n2164) );
  or2 U2308 ( .A1(n2165), .A2(n2164), .Z(n2166) );
  and2 U2309 ( .A1(n2944), .A2(n2166), .Z(n1461) );
  inv1 U2310 ( .I(n2166), .ZN(n2167) );
  and2 U2311 ( .A1(n2168), .A2(n2167), .Z(n1462) );
  inv1 U2312 ( .I(k5), .ZN(n3698) );
  inv1 U2313 ( .I(m5), .ZN(n3697) );
  inv1 U2314 ( .I(c6), .ZN(n3687) );
  inv1 U2315 ( .I(a6), .ZN(n3689) );
  inv1 U2316 ( .I(z5), .ZN(n3690) );
  inv1 U2317 ( .I(w5), .ZN(n3693) );
  inv1 U2318 ( .I(b6), .ZN(n3688) );
  inv1 U2319 ( .I(y5), .ZN(n3691) );
  inv1 U2320 ( .I(w6), .ZN(n3686) );
  or2 U2321 ( .A1(n1947), .A2(n1292), .Z(n2251) );
  and2 U2322 ( .A1(n2169), .A2(f), .Z(n2171) );
  and2 U2323 ( .A1(m0), .A2(n1928), .Z(n2170) );
  or2 U2324 ( .A1(n2171), .A2(n2170), .Z(n2398) );
  and2 U2325 ( .A1(n2251), .A2(n2398), .Z(n1152) );
  and2 U2326 ( .A1(n2172), .A2(f), .Z(n2174) );
  and2 U2327 ( .A1(x), .A2(n2122), .Z(n2173) );
  or2 U2328 ( .A1(n2174), .A2(n2173), .Z(n715) );
  or2 U2329 ( .A1(n1962), .A2(n1310), .Z(n2234) );
  or2 U2330 ( .A1(n2234), .A2(n715), .Z(n1153) );
  and2 U2331 ( .A1(n715), .A2(n2234), .Z(n1151) );
  inv1 U2332 ( .I(v6), .ZN(n2175) );
  and2 U2333 ( .A1(n2175), .A2(f), .Z(n2177) );
  and2 U2334 ( .A1(y), .A2(n2116), .Z(n2176) );
  or2 U2335 ( .A1(n2177), .A2(n2176), .Z(n719) );
  or2 U2336 ( .A1(n1952), .A2(n1305), .Z(n2833) );
  or2 U2337 ( .A1(n2833), .A2(n719), .Z(n1148) );
  inv1 U2338 ( .I(x5), .ZN(n3692) );
  inv1 U2339 ( .I(p5), .ZN(n3694) );
  inv1 U2340 ( .I(o5), .ZN(n3695) );
  inv1 U2341 ( .I(b1), .ZN(n3699) );
  inv1 U2342 ( .I(n5), .ZN(n3696) );
  and2 U2343 ( .A1(g1), .A2(n2072), .Z(n2178) );
  or2 U2344 ( .A1(n2178), .A2(n1350), .Z(n812) );
  and2 U2345 ( .A1(e1), .A2(n2120), .Z(n2179) );
  or2 U2346 ( .A1(n2179), .A2(n1078), .Z(n803) );
  and2 U2347 ( .A1(n812), .A2(n2101), .Z(n2182) );
  inv1 U2348 ( .I(o2), .ZN(n2180) );
  and2 U2349 ( .A1(n2180), .A2(f), .Z(n2181) );
  or2 U2350 ( .A1(n2181), .A2(n2104), .Z(n2301) );
  inv1 U2351 ( .I(n2301), .ZN(n2303) );
  or2 U2352 ( .A1(n2303), .A2(n803), .Z(n2883) );
  and2 U2353 ( .A1(n2182), .A2(n2883), .Z(n1069) );
  and2 U2354 ( .A1(n803), .A2(n2303), .Z(n1070) );
  and2 U2355 ( .A1(u0), .A2(n1944), .Z(n2183) );
  or2 U2356 ( .A1(n2183), .A2(n1081), .Z(n836) );
  inv1 U2357 ( .I(n2), .ZN(n2184) );
  and2 U2358 ( .A1(n2184), .A2(f), .Z(n2185) );
  or2 U2359 ( .A1(n2185), .A2(n2104), .Z(n2302) );
  inv1 U2360 ( .I(n2302), .ZN(n2300) );
  or2 U2361 ( .A1(n2300), .A2(n836), .Z(n1067) );
  and2 U2362 ( .A1(n836), .A2(n2300), .Z(n1066) );
  and2 U2363 ( .A1(f1), .A2(n2118), .Z(n2186) );
  or2 U2364 ( .A1(n2186), .A2(n1086), .Z(n841) );
  inv1 U2365 ( .I(m2), .ZN(n2187) );
  and2 U2366 ( .A1(n2187), .A2(f), .Z(n2188) );
  or2 U2367 ( .A1(n2188), .A2(n3708), .Z(n2299) );
  inv1 U2368 ( .I(n2299), .ZN(n2908) );
  or2 U2369 ( .A1(n2908), .A2(n841), .Z(n1063) );
  or2 U2370 ( .A1(n1943), .A2(n1138), .Z(n2192) );
  inv1 U2371 ( .I(n2192), .ZN(n2851) );
  inv1 U2372 ( .I(w2), .ZN(n2189) );
  and2 U2373 ( .A1(n2189), .A2(f), .Z(n2190) );
  or2 U2374 ( .A1(n2190), .A2(n2104), .Z(n2857) );
  and2 U2375 ( .A1(n2851), .A2(n2857), .Z(n1043) );
  inv1 U2376 ( .I(n2857), .ZN(n2191) );
  and2 U2377 ( .A1(n2192), .A2(n2191), .Z(n1044) );
  inv1 U2378 ( .I(s2), .ZN(n2193) );
  and2 U2379 ( .A1(n2193), .A2(f), .Z(n2194) );
  or2 U2380 ( .A1(n2194), .A2(n2104), .Z(n2726) );
  inv1 U2381 ( .I(n2726), .ZN(n2873) );
  or2 U2382 ( .A1(n1941), .A2(n1336), .Z(n2197) );
  inv1 U2383 ( .I(t2), .ZN(n2195) );
  and2 U2384 ( .A1(n2195), .A2(f), .Z(n2196) );
  or2 U2385 ( .A1(n2196), .A2(n2104), .Z(n2870) );
  inv1 U2386 ( .I(n2870), .ZN(n2867) );
  and2 U2387 ( .A1(n2197), .A2(n2867), .Z(n2199) );
  inv1 U2388 ( .I(n2197), .ZN(n2848) );
  and2 U2389 ( .A1(n2848), .A2(n2870), .Z(n2198) );
  or2 U2390 ( .A1(n2199), .A2(n2198), .Z(n2201) );
  inv1 U2391 ( .I(n2201), .ZN(n2200) );
  and2 U2392 ( .A1(n2873), .A2(n2200), .Z(n1033) );
  and2 U2393 ( .A1(n2726), .A2(n2201), .Z(n1034) );
  inv1 U2394 ( .I(v2), .ZN(n2202) );
  and2 U2395 ( .A1(n2202), .A2(f), .Z(n2203) );
  or2 U2396 ( .A1(n2203), .A2(n3709), .Z(n2860) );
  inv1 U2397 ( .I(n2860), .ZN(n2206) );
  inv1 U2398 ( .I(u2), .ZN(n2204) );
  and2 U2399 ( .A1(n2204), .A2(f), .Z(n2205) );
  or2 U2400 ( .A1(n2205), .A2(n2104), .Z(n2861) );
  and2 U2401 ( .A1(n2206), .A2(n2861), .Z(n1016) );
  inv1 U2402 ( .I(n2861), .ZN(n2207) );
  and2 U2403 ( .A1(n2860), .A2(n2207), .Z(n1017) );
  and2 U2404 ( .A1(q2), .A2(f), .Z(n2208) );
  and2 U2407 ( .A1(s1), .A2(n2889), .Z(n2211) );
  inv1 U2408 ( .I(s1), .ZN(n2209) );
  and2 U2409 ( .A1(n2209), .A2(n2213), .Z(n2210) );
  or2 U2410 ( .A1(n2211), .A2(n2210), .Z(n2212) );
  and2 U2411 ( .A1(n2111), .A2(n2212), .Z(n2219) );
  and2 U2412 ( .A1(a3), .A2(n2889), .Z(n2216) );
  inv1 U2413 ( .I(a3), .ZN(n2214) );
  and2 U2414 ( .A1(n2214), .A2(n2213), .Z(n2215) );
  and2 U2416 ( .A1(f), .A2(n2217), .Z(n2218) );
  or2 U2417 ( .A1(n2219), .A2(n2218), .Z(n1015) );
  and2 U2419 ( .A1(z2), .A2(f), .Z(n2222) );
  inv1 U2420 ( .I(r1), .ZN(n2220) );
  or2 U2421 ( .A1(n2080), .A2(n2220), .Z(n2221) );
  inv1 U2422 ( .I(n2221), .ZN(n2457) );
  and2 U2424 ( .A1(n2223), .A2(n2224), .Z(n2226) );
  or2 U2428 ( .A1(n1931), .A2(n1182), .Z(n2228) );
  inv1 U2429 ( .I(n2228), .ZN(n2749) );
  or2 U2430 ( .A1(n1935), .A2(n1184), .Z(n2227) );
  and2 U2431 ( .A1(n2749), .A2(n2227), .Z(n990) );
  inv1 U2432 ( .I(n2227), .ZN(n2745) );
  and2 U2433 ( .A1(n2228), .A2(n2745), .Z(n991) );
  inv1 U2434 ( .I(n2833), .ZN(n2229) );
  or2 U2435 ( .A1(n1933), .A2(n1300), .Z(n2832) );
  and2 U2436 ( .A1(n2229), .A2(n2832), .Z(n2232) );
  inv1 U2437 ( .I(n2832), .ZN(n2230) );
  and2 U2438 ( .A1(n2833), .A2(n2230), .Z(n2231) );
  or2 U2439 ( .A1(n2232), .A2(n2231), .Z(n2233) );
  or2 U2440 ( .A1(n2233), .A2(n2234), .Z(n979) );
  inv1 U2441 ( .I(n2233), .ZN(n2236) );
  inv1 U2442 ( .I(n2234), .ZN(n2235) );
  or2 U2443 ( .A1(n2236), .A2(n2235), .Z(n3704) );
  inv1 U2446 ( .I(n2242), .ZN(n2817) );
  inv1 U2448 ( .I(i1), .ZN(n2238) );
  and2 U2449 ( .A1(n2238), .A2(n2242), .Z(n2239) );
  or2 U2450 ( .A1(n2240), .A2(n2239), .Z(n2241) );
  and2 U2451 ( .A1(n2072), .A2(n2241), .Z(n2248) );
  and2 U2452 ( .A1(q3), .A2(n2817), .Z(n2245) );
  inv1 U2453 ( .I(q3), .ZN(n2243) );
  and2 U2454 ( .A1(n2243), .A2(n2242), .Z(n2244) );
  or2 U2455 ( .A1(n2245), .A2(n2244), .Z(n2246) );
  inv1 U2458 ( .I(n2251), .ZN(n2730) );
  and2 U2459 ( .A1(p3), .A2(f), .Z(n2249) );
  or2 U2460 ( .A1(n2249), .A2(n1948), .Z(n2250) );
  and2 U2461 ( .A1(n2730), .A2(n2250), .Z(n2253) );
  inv1 U2462 ( .I(n2250), .ZN(n2735) );
  and2 U2463 ( .A1(n2251), .A2(n2735), .Z(n2252) );
  or2 U2464 ( .A1(n2253), .A2(n2252), .Z(n959) );
  or2 U2465 ( .A1(n1937), .A2(n1189), .Z(n2733) );
  or2 U2466 ( .A1(n2733), .A2(n950), .Z(n947) );
  inv1 U2469 ( .I(b4), .ZN(n2258) );
  inv1 U2471 ( .I(m), .ZN(n2255) );
  or2 U2472 ( .A1(f), .A2(n2255), .Z(n2256) );
  inv1 U2473 ( .I(n2256), .ZN(n2535) );
  and2 U2475 ( .A1(n2258), .A2(n2261), .Z(n2260) );
  or2 U2478 ( .A1(n2260), .A2(n2259), .Z(n915) );
  and2 U2479 ( .A1(n439), .A2(n2261), .Z(n2263) );
  and2 U2480 ( .A1(n), .A2(n2793), .Z(n2262) );
  or2 U2481 ( .A1(n2263), .A2(n2262), .Z(n2264) );
  and2 U2482 ( .A1(n2120), .A2(n2264), .Z(n2265) );
  or2 U2483 ( .A1(n2265), .A2(n914), .Z(n904) );
  and2 U2484 ( .A1(x3), .A2(f), .Z(n2266) );
  or2 U2485 ( .A1(n2266), .A2(n1927), .Z(n2268) );
  and2 U2486 ( .A1(w3), .A2(f), .Z(n2267) );
  or2 U2487 ( .A1(n2267), .A2(n1924), .Z(n2269) );
  inv1 U2488 ( .I(n2269), .ZN(n2807) );
  and2 U2489 ( .A1(n2268), .A2(n2807), .Z(n2271) );
  inv1 U2490 ( .I(n2268), .ZN(n2761) );
  and2 U2491 ( .A1(n2761), .A2(n2269), .Z(n2270) );
  or2 U2492 ( .A1(n2271), .A2(n2270), .Z(n903) );
  and2 U2493 ( .A1(v3), .A2(f), .Z(n2272) );
  or2 U2494 ( .A1(n1945), .A2(n2272), .Z(n2274) );
  and2 U2495 ( .A1(u3), .A2(f), .Z(n2273) );
  or2 U2496 ( .A1(n2273), .A2(n1950), .Z(n2275) );
  inv1 U2497 ( .I(n2275), .ZN(n2779) );
  and2 U2498 ( .A1(n2274), .A2(n2779), .Z(n2277) );
  inv1 U2499 ( .I(n2274), .ZN(n2771) );
  and2 U2500 ( .A1(n2771), .A2(n2275), .Z(n2276) );
  or2 U2501 ( .A1(n2277), .A2(n2276), .Z(n2278) );
  or2 U2502 ( .A1(n1939), .A2(n1279), .Z(n2765) );
  inv1 U2503 ( .I(n2765), .ZN(n2775) );
  and2 U2504 ( .A1(n2278), .A2(n2775), .Z(n2281) );
  inv1 U2505 ( .I(n2278), .ZN(n2279) );
  and2 U2506 ( .A1(n2279), .A2(n2765), .Z(n2280) );
  or2 U2507 ( .A1(n2281), .A2(n2280), .Z(n2282) );
  inv1 U2508 ( .I(n2282), .ZN(n3679) );
  and2 U2510 ( .A1(a4), .A2(f), .Z(n2283) );
  or2 U2511 ( .A1(n2283), .A2(n1949), .Z(n2285) );
  and2 U2512 ( .A1(y3), .A2(f), .Z(n2284) );
  or2 U2513 ( .A1(n2284), .A2(n1929), .Z(n2286) );
  inv1 U2514 ( .I(n2286), .ZN(n2784) );
  and2 U2515 ( .A1(n2285), .A2(n2784), .Z(n2288) );
  inv1 U2516 ( .I(n2285), .ZN(n2790) );
  and2 U2517 ( .A1(n2790), .A2(n2286), .Z(n2287) );
  or2 U2518 ( .A1(n2288), .A2(n2287), .Z(n889) );
  inv1 U2519 ( .I(n893), .ZN(n2292) );
  and2 U2520 ( .A1(z3), .A2(f), .Z(n2291) );
  inv1 U2521 ( .I(h), .ZN(n2289) );
  or2 U2522 ( .A1(f), .A2(n2289), .Z(n2290) );
  inv1 U2523 ( .I(n2290), .ZN(n2568) );
  or2 U2524 ( .A1(n2291), .A2(n2568), .Z(n2293) );
  inv1 U2526 ( .I(n2293), .ZN(n2786) );
  and2 U2527 ( .A1(n893), .A2(n2786), .Z(n2294) );
  inv1 U2529 ( .I(l2), .ZN(n2296) );
  and2 U2530 ( .A1(n2296), .A2(f), .Z(n2297) );
  or2 U2531 ( .A1(n2297), .A2(n2104), .Z(n2298) );
  or2 U2532 ( .A1(n2298), .A2(n2908), .Z(n3702) );
  inv1 U2533 ( .I(n2298), .ZN(n2907) );
  or2 U2534 ( .A1(n2907), .A2(n2299), .Z(n880) );
  and2 U2535 ( .A1(n2301), .A2(n2300), .Z(n873) );
  and2 U2536 ( .A1(n2303), .A2(n2302), .Z(n874) );
  and2 U2537 ( .A1(k2), .A2(f), .Z(n2309) );
  inv1 U2538 ( .I(j2), .ZN(n2304) );
  and2 U2539 ( .A1(n2304), .A2(p2), .Z(n2307) );
  inv1 U2540 ( .I(p2), .ZN(n2305) );
  and2 U2541 ( .A1(j2), .A2(n2305), .Z(n2306) );
  or2 U2542 ( .A1(n2307), .A2(n2306), .Z(n2310) );
  and2 U2543 ( .A1(n2101), .A2(n2310), .Z(n2308) );
  and2 U2544 ( .A1(n2309), .A2(n2308), .Z(n855) );
  and2 U2545 ( .A1(f), .A2(n2101), .Z(n2314) );
  inv1 U2546 ( .I(k2), .ZN(n2312) );
  inv1 U2547 ( .I(n2310), .ZN(n2311) );
  and2 U2548 ( .A1(n2312), .A2(n2311), .Z(n2313) );
  and2 U2549 ( .A1(n2314), .A2(n2313), .Z(n856) );
  and2 U2550 ( .A1(v0), .A2(n1946), .Z(n2315) );
  or2 U2551 ( .A1(n2315), .A2(n1090), .Z(n840) );
  inv1 U2552 ( .I(n840), .ZN(n3678) );
  inv1 U2553 ( .I(n841), .ZN(n3680) );
  inv1 U2554 ( .I(q5), .ZN(n2316) );
  and2 U2555 ( .A1(n2316), .A2(f), .Z(n2318) );
  inv1 U2556 ( .I(n829), .ZN(n2317) );
  or2 U2557 ( .A1(n2318), .A2(n2317), .Z(n3701) );
  inv1 U2558 ( .I(n3701), .ZN(n827) );
  inv1 U2559 ( .I(n816), .ZN(n815) );
  inv1 U2560 ( .I(n803), .ZN(n3681) );
  and2 U2561 ( .A1(n813), .A2(n2116), .Z(n2319) );
  or2 U2562 ( .A1(n2319), .A2(n807), .Z(n804) );
  inv1 U2563 ( .I(n804), .ZN(n802) );
  and2 U2564 ( .A1(n824), .A2(n1930), .Z(n2320) );
  or2 U2565 ( .A1(n2320), .A2(n818), .Z(n798) );
  inv1 U2566 ( .I(d6), .ZN(n2321) );
  and2 U2568 ( .A1(e0), .A2(n3710), .Z(n2322) );
  and2 U2571 ( .A1(f0), .A2(n3677), .Z(n2325) );
  inv1 U2572 ( .I(f0), .ZN(n2792) );
  and2 U2573 ( .A1(n2792), .A2(n767), .Z(n2324) );
  or2 U2574 ( .A1(n2325), .A2(n2324), .Z(n2326) );
  and2 U2575 ( .A1(n1930), .A2(n2326), .Z(n2327) );
  or2 U2576 ( .A1(n2327), .A2(n761), .Z(n2328) );
  inv1 U2577 ( .I(n2328), .ZN(n3676) );
  inv1 U2578 ( .I(j6), .ZN(n2617) );
  and2 U2579 ( .A1(n2617), .A2(f), .Z(n2330) );
  and2 U2580 ( .A1(q), .A2(n1951), .Z(n2329) );
  or2 U2581 ( .A1(n2330), .A2(n2329), .Z(n2334) );
  inv1 U2582 ( .I(i6), .ZN(n2331) );
  and2 U2583 ( .A1(n2331), .A2(f), .Z(n2333) );
  and2 U2584 ( .A1(g0), .A2(n2118), .Z(n2332) );
  or2 U2585 ( .A1(n2333), .A2(n2332), .Z(n2335) );
  inv1 U2586 ( .I(n2335), .ZN(n2762) );
  and2 U2587 ( .A1(n2334), .A2(n2762), .Z(n2337) );
  inv1 U2588 ( .I(n2334), .ZN(n2806) );
  and2 U2589 ( .A1(n2806), .A2(n2335), .Z(n2336) );
  or2 U2590 ( .A1(n2337), .A2(n2336), .Z(n2338) );
  inv1 U2591 ( .I(n2338), .ZN(n3675) );
  inv1 U2592 ( .I(l6), .ZN(n2339) );
  and2 U2593 ( .A1(n2339), .A2(f), .Z(n2341) );
  and2 U2594 ( .A1(s), .A2(n1930), .Z(n2340) );
  inv1 U2596 ( .I(m6), .ZN(n2342) );
  and2 U2597 ( .A1(n2342), .A2(f), .Z(n2344) );
  and2 U2598 ( .A1(t), .A2(n2111), .Z(n2343) );
  or2 U2599 ( .A1(n2344), .A2(n2343), .Z(n2766) );
  inv1 U2600 ( .I(k6), .ZN(n2345) );
  and2 U2601 ( .A1(n2345), .A2(f), .Z(n2347) );
  and2 U2602 ( .A1(r), .A2(n2122), .Z(n2346) );
  or2 U2603 ( .A1(n2347), .A2(n2346), .Z(n2348) );
  inv1 U2604 ( .I(n2348), .ZN(n2770) );
  and2 U2605 ( .A1(n2766), .A2(n2770), .Z(n2350) );
  inv1 U2606 ( .I(n2766), .ZN(n2776) );
  and2 U2607 ( .A1(n2776), .A2(n2348), .Z(n2349) );
  or2 U2608 ( .A1(n2350), .A2(n2349), .Z(n2353) );
  inv1 U2609 ( .I(n2353), .ZN(n2351) );
  and2 U2610 ( .A1(n2352), .A2(n2351), .Z(n2355) );
  inv1 U2611 ( .I(n2352), .ZN(n2780) );
  and2 U2612 ( .A1(n2780), .A2(n2353), .Z(n2354) );
  or2 U2613 ( .A1(n2355), .A2(n2354), .Z(n744) );
  inv1 U2614 ( .I(n745), .ZN(n740) );
  inv1 U2615 ( .I(h6), .ZN(n2356) );
  and2 U2616 ( .A1(n2356), .A2(f), .Z(n2358) );
  and2 U2617 ( .A1(i0), .A2(n1930), .Z(n2357) );
  or2 U2618 ( .A1(n2358), .A2(n2357), .Z(n2362) );
  inv1 U2619 ( .I(f6), .ZN(n2359) );
  and2 U2620 ( .A1(n2359), .A2(f), .Z(n2361) );
  and2 U2621 ( .A1(h0), .A2(n2122), .Z(n2360) );
  or2 U2622 ( .A1(n2361), .A2(n2360), .Z(n2363) );
  inv1 U2623 ( .I(n2363), .ZN(n2791) );
  and2 U2624 ( .A1(n2362), .A2(n2791), .Z(n2365) );
  inv1 U2625 ( .I(n2362), .ZN(n2785) );
  and2 U2626 ( .A1(n2785), .A2(n2363), .Z(n2364) );
  or2 U2627 ( .A1(n2365), .A2(n2364), .Z(n2366) );
  inv1 U2628 ( .I(n2366), .ZN(n3674) );
  and2 U2629 ( .A1(n2018), .A2(f), .Z(n2368) );
  and2 U2630 ( .A1(j0), .A2(n1944), .Z(n2367) );
  or2 U2631 ( .A1(n2368), .A2(n2367), .Z(n2369) );
  inv1 U2632 ( .I(n2369), .ZN(n2787) );
  and2 U2633 ( .A1(n737), .A2(n2787), .Z(n2372) );
  inv1 U2634 ( .I(n737), .ZN(n2370) );
  inv1 U2638 ( .I(s6), .ZN(n2374) );
  and2 U2639 ( .A1(n2374), .A2(f), .Z(n2376) );
  and2 U2640 ( .A1(n0), .A2(n1930), .Z(n2375) );
  or2 U2641 ( .A1(n2376), .A2(n2375), .Z(n725) );
  inv1 U2642 ( .I(n725), .ZN(n3672) );
  inv1 U2643 ( .I(r6), .ZN(n2377) );
  and2 U2644 ( .A1(n2377), .A2(f), .Z(n2379) );
  and2 U2645 ( .A1(o0), .A2(n1946), .Z(n2378) );
  or2 U2646 ( .A1(n2379), .A2(n2378), .Z(n726) );
  inv1 U2647 ( .I(n726), .ZN(n3671) );
  and2 U2648 ( .A1(z), .A2(n1944), .Z(n2380) );
  or2 U2649 ( .A1(n2380), .A2(n1297), .Z(n2831) );
  inv1 U2650 ( .I(n2831), .ZN(n3670) );
  inv1 U2651 ( .I(o6), .ZN(n2621) );
  and2 U2652 ( .A1(n2621), .A2(f), .Z(n2382) );
  and2 U2653 ( .A1(k0), .A2(n2072), .Z(n2381) );
  or2 U2654 ( .A1(n2382), .A2(n2381), .Z(n2389) );
  inv1 U2655 ( .I(n2389), .ZN(n2816) );
  and2 U2656 ( .A1(v), .A2(n2816), .Z(n2385) );
  inv1 U2657 ( .I(v), .ZN(n2383) );
  and2 U2658 ( .A1(n2383), .A2(n2389), .Z(n2384) );
  or2 U2659 ( .A1(n2385), .A2(n2384), .Z(n2386) );
  and2 U2660 ( .A1(n2049), .A2(n2386), .Z(n2393) );
  or2 U2661 ( .A1(n2816), .A2(n6), .Z(n2387) );
  and2 U2662 ( .A1(f), .A2(n2387), .Z(n2391) );
  inv1 U2663 ( .I(n6), .ZN(n2388) );
  or2 U2664 ( .A1(n2389), .A2(n2388), .Z(n2390) );
  and2 U2665 ( .A1(n2391), .A2(n2390), .Z(n2392) );
  or2 U2666 ( .A1(n2393), .A2(n2392), .Z(n692) );
  inv1 U2667 ( .I(n2398), .ZN(n2729) );
  inv1 U2668 ( .I(p6), .ZN(n2394) );
  and2 U2669 ( .A1(n2394), .A2(f), .Z(n2396) );
  and2 U2670 ( .A1(l0), .A2(n2118), .Z(n2395) );
  or2 U2671 ( .A1(n2396), .A2(n2395), .Z(n2397) );
  and2 U2672 ( .A1(n2729), .A2(n2397), .Z(n2400) );
  inv1 U2673 ( .I(n2397), .ZN(n2734) );
  and2 U2674 ( .A1(n2398), .A2(n2734), .Z(n2399) );
  or2 U2675 ( .A1(n2400), .A2(n2399), .Z(n691) );
  inv1 U2676 ( .I(q6), .ZN(n2401) );
  and2 U2677 ( .A1(n2401), .A2(f), .Z(n2403) );
  and2 U2678 ( .A1(w), .A2(n1944), .Z(n2402) );
  or2 U2679 ( .A1(n2403), .A2(n2402), .Z(n683) );
  and2 U2680 ( .A1(s0), .A2(n2049), .Z(n2404) );
  or2 U2681 ( .A1(n2404), .A2(n1135), .Z(n671) );
  inv1 U2682 ( .I(n671), .ZN(n3669) );
  and2 U2683 ( .A1(b0), .A2(n1930), .Z(n2405) );
  or2 U2684 ( .A1(n2405), .A2(n1317), .Z(n672) );
  inv1 U2685 ( .I(n672), .ZN(n3668) );
  and2 U2686 ( .A1(r0), .A2(n1930), .Z(n2406) );
  or2 U2687 ( .A1(n2406), .A2(n1333), .Z(n665) );
  inv1 U2688 ( .I(n665), .ZN(n3667) );
  and2 U2689 ( .A1(c1), .A2(n2120), .Z(n2407) );
  or2 U2690 ( .A1(n2407), .A2(n1328), .Z(n666) );
  inv1 U2691 ( .I(n666), .ZN(n3666) );
  and2 U2692 ( .A1(d1), .A2(n3710), .Z(n2408) );
  or2 U2693 ( .A1(n2408), .A2(n1345), .Z(n660) );
  and2 U2694 ( .A1(a0), .A2(n1951), .Z(n2409) );
  or2 U2695 ( .A1(n2409), .A2(n1338), .Z(n643) );
  inv1 U2696 ( .I(n643), .ZN(n3665) );
  and2 U2697 ( .A1(t0), .A2(n2119), .Z(n2410) );
  or2 U2698 ( .A1(n2410), .A2(n1341), .Z(n644) );
  inv1 U2699 ( .I(n644), .ZN(n3664) );
  inv1 U2700 ( .I(u5), .ZN(n2633) );
  and2 U2702 ( .A1(c0), .A2(n2119), .Z(n2411) );
  and2 U2705 ( .A1(p0), .A2(n2888), .Z(n2415) );
  inv1 U2706 ( .I(p0), .ZN(n2413) );
  and2 U2707 ( .A1(n2413), .A2(n2419), .Z(n2414) );
  or2 U2708 ( .A1(n2415), .A2(n2414), .Z(n2416) );
  and2 U2709 ( .A1(n2119), .A2(n2416), .Z(n2423) );
  and2 U2711 ( .A1(f), .A2(n2417), .Z(n2421) );
  inv1 U2712 ( .I(t5), .ZN(n2418) );
  or2 U2713 ( .A1(n2419), .A2(n2418), .Z(n2420) );
  and2 U2714 ( .A1(n2421), .A2(n2420), .Z(n2422) );
  or2 U2715 ( .A1(n2423), .A2(n2422), .Z(n639) );
  inv1 U2716 ( .I(n628), .ZN(n2426) );
  inv1 U2717 ( .I(v5), .ZN(n2636) );
  and2 U2718 ( .A1(n2636), .A2(f), .Z(n2425) );
  and2 U2719 ( .A1(q0), .A2(n2120), .Z(n2424) );
  or2 U2720 ( .A1(n2425), .A2(n2424), .Z(n2427) );
  and2 U2721 ( .A1(n2426), .A2(n2427), .Z(n2429) );
  inv1 U2722 ( .I(n2427), .ZN(n2841) );
  and2 U2723 ( .A1(n628), .A2(n2841), .Z(n2428) );
  inv1 U2725 ( .I(b2), .ZN(n2430) );
  and2 U2726 ( .A1(n2430), .A2(f), .Z(n2431) );
  inv1 U2728 ( .I(n2579), .ZN(n2578) );
  inv1 U2729 ( .I(c2), .ZN(n2432) );
  and2 U2732 ( .A1(n2578), .A2(n2627), .Z(n574) );
  inv1 U2733 ( .I(n2627), .ZN(n2651) );
  and2 U2734 ( .A1(n2579), .A2(n2651), .Z(n575) );
  and2 U2735 ( .A1(w1), .A2(n2107), .Z(n2434) );
  or2 U2736 ( .A1(n2434), .A2(n1921), .Z(n2634) );
  inv1 U2737 ( .I(n2015), .ZN(n2635) );
  and2 U2738 ( .A1(g2), .A2(f), .Z(n2436) );
  and2 U2739 ( .A1(s1), .A2(n2120), .Z(n2435) );
  or2 U2740 ( .A1(n2436), .A2(n2435), .Z(n2437) );
  and2 U2741 ( .A1(n2635), .A2(n2437), .Z(n2443) );
  inv1 U2742 ( .I(g2), .ZN(n2438) );
  and2 U2743 ( .A1(n2438), .A2(f), .Z(n2440) );
  and2 U2744 ( .A1(n2209), .A2(n2120), .Z(n2439) );
  or2 U2745 ( .A1(n2440), .A2(n2439), .Z(n2441) );
  and2 U2746 ( .A1(n2634), .A2(n2441), .Z(n2442) );
  or2 U2747 ( .A1(n2443), .A2(n2442), .Z(n572) );
  inv1 U2748 ( .I(a2), .ZN(n2444) );
  inv1 U2751 ( .I(y1), .ZN(n2446) );
  and2 U2752 ( .A1(n2446), .A2(f), .Z(n2447) );
  inv1 U2754 ( .I(z1), .ZN(n2448) );
  and2 U2755 ( .A1(n2448), .A2(f), .Z(n2449) );
  or2 U2756 ( .A1(n2449), .A2(n3707), .Z(n2576) );
  inv1 U2757 ( .I(n2576), .ZN(n2450) );
  and2 U2760 ( .A1(n2675), .A2(n2576), .Z(n2451) );
  or2 U2761 ( .A1(n2452), .A2(n2451), .Z(n2454) );
  inv1 U2762 ( .I(n2454), .ZN(n2453) );
  and2 U2763 ( .A1(n2678), .A2(n2453), .Z(n2456) );
  inv1 U2764 ( .I(n2678), .ZN(n2689) );
  and2 U2765 ( .A1(n2689), .A2(n2454), .Z(n2455) );
  or2 U2766 ( .A1(n2456), .A2(n2455), .Z(n568) );
  inv1 U2767 ( .I(n566), .ZN(n565) );
  and2 U2768 ( .A1(f2), .A2(n2079), .Z(n2458) );
  and2 U2769 ( .A1(d2), .A2(f), .Z(n2459) );
  or2 U2770 ( .A1(n2459), .A2(n1943), .Z(n2460) );
  inv1 U2771 ( .I(n2460), .ZN(n2630) );
  and2 U2772 ( .A1(n2637), .A2(n2630), .Z(n2462) );
  and2 U2773 ( .A1(n1965), .A2(n2460), .Z(n2461) );
  or2 U2774 ( .A1(n2462), .A2(n2461), .Z(n557) );
  and2 U2775 ( .A1(e2), .A2(f), .Z(n2463) );
  or2 U2776 ( .A1(n2463), .A2(n1941), .Z(n2464) );
  inv1 U2777 ( .I(n2464), .ZN(n2640) );
  and2 U2778 ( .A1(n560), .A2(n2640), .Z(n2467) );
  inv1 U2779 ( .I(n560), .ZN(n2465) );
  and2 U2780 ( .A1(n2465), .A2(n2464), .Z(n2466) );
  or2 U2781 ( .A1(n2467), .A2(n2466), .Z(n2468) );
  inv1 U2783 ( .I(g4), .ZN(n2469) );
  and2 U2784 ( .A1(n2469), .A2(f), .Z(n2470) );
  or2 U2785 ( .A1(n2470), .A2(n3708), .Z(n2586) );
  inv1 U2786 ( .I(i4), .ZN(n2471) );
  and2 U2787 ( .A1(n2471), .A2(n2107), .Z(n2472) );
  inv1 U2789 ( .I(n2594), .ZN(n2473) );
  and2 U2790 ( .A1(n2586), .A2(n2473), .Z(n2475) );
  inv1 U2791 ( .I(n2586), .ZN(n2702) );
  and2 U2792 ( .A1(n2702), .A2(n2594), .Z(n2474) );
  or2 U2793 ( .A1(n2475), .A2(n2474), .Z(n2476) );
  inv1 U2794 ( .I(n2476), .ZN(n3662) );
  inv1 U2795 ( .I(c4), .ZN(n2477) );
  and2 U2796 ( .A1(n2477), .A2(f), .Z(n2478) );
  inv1 U2798 ( .I(j4), .ZN(n2479) );
  and2 U2799 ( .A1(n2479), .A2(n2080), .Z(n2480) );
  inv1 U2801 ( .I(n2591), .ZN(n2703) );
  and2 U2802 ( .A1(n2590), .A2(n2703), .Z(n2482) );
  inv1 U2803 ( .I(n2590), .ZN(n2589) );
  and2 U2804 ( .A1(n2589), .A2(n1992), .Z(n2481) );
  or2 U2805 ( .A1(n2482), .A2(n2481), .Z(n538) );
  inv1 U2806 ( .I(h4), .ZN(n2483) );
  and2 U2807 ( .A1(n2483), .A2(f), .Z(n2484) );
  or2 U2808 ( .A1(n2484), .A2(n2104), .Z(n2597) );
  inv1 U2809 ( .I(n2597), .ZN(n2485) );
  or2 U2810 ( .A1(n2485), .A2(n3707), .Z(n2495) );
  inv1 U2811 ( .I(n2495), .ZN(n2492) );
  or2 U2812 ( .A1(n1951), .A2(e4), .Z(n2487) );
  inv1 U2813 ( .I(n2487), .ZN(n2486) );
  and2 U2814 ( .A1(n529), .A2(n2486), .Z(n2491) );
  inv1 U2815 ( .I(n529), .ZN(n2488) );
  and2 U2816 ( .A1(n2488), .A2(n2487), .Z(n2489) );
  or2 U2817 ( .A1(n2489), .A2(n2104), .Z(n2490) );
  or2 U2818 ( .A1(n2491), .A2(n2490), .Z(n2493) );
  and2 U2819 ( .A1(n2492), .A2(n2493), .Z(n519) );
  inv1 U2820 ( .I(n2493), .ZN(n2494) );
  and2 U2821 ( .A1(n2495), .A2(n2494), .Z(n520) );
  and2 U2822 ( .A1(k4), .A2(f), .Z(n2496) );
  or2 U2823 ( .A1(n2496), .A2(n1925), .Z(n2622) );
  inv1 U2824 ( .I(n2622), .ZN(n2608) );
  and2 U2825 ( .A1(u4), .A2(f), .Z(n2498) );
  and2 U2826 ( .A1(i1), .A2(n1930), .Z(n2497) );
  or2 U2827 ( .A1(n2498), .A2(n2497), .Z(n2499) );
  and2 U2828 ( .A1(n2608), .A2(n2499), .Z(n2505) );
  inv1 U2829 ( .I(u4), .ZN(n2500) );
  and2 U2830 ( .A1(n2500), .A2(f), .Z(n2502) );
  and2 U2831 ( .A1(n2238), .A2(n1930), .Z(n2501) );
  or2 U2832 ( .A1(n2502), .A2(n2501), .Z(n2503) );
  and2 U2833 ( .A1(n1909), .A2(n2503), .Z(n2504) );
  or2 U2834 ( .A1(n2505), .A2(n2504), .Z(n475) );
  and2 U2835 ( .A1(q4), .A2(f), .Z(n2506) );
  or2 U2836 ( .A1(n2506), .A2(n1931), .Z(n2508) );
  inv1 U2837 ( .I(n2508), .ZN(n2673) );
  and2 U2838 ( .A1(n2507), .A2(n2673), .Z(n2511) );
  and2 U2839 ( .A1(n2509), .A2(n2508), .Z(n2510) );
  or2 U2840 ( .A1(n2511), .A2(n2510), .Z(n474) );
  and2 U2841 ( .A1(n1985), .A2(n2512), .Z(n2516) );
  and2 U2842 ( .A1(n2514), .A2(n2513), .Z(n2515) );
  or2 U2843 ( .A1(n2516), .A2(n2515), .Z(n2519) );
  inv1 U2844 ( .I(n2519), .ZN(n2517) );
  and2 U2845 ( .A1(n2518), .A2(n2517), .Z(n2522) );
  and2 U2846 ( .A1(n2520), .A2(n2519), .Z(n2521) );
  or2 U2847 ( .A1(n2522), .A2(n2521), .Z(n471) );
  inv1 U2848 ( .I(n469), .ZN(n468) );
  or2 U2850 ( .A1(n2523), .A2(n1948), .Z(n2525) );
  and2 U2851 ( .A1(r4), .A2(f), .Z(n2524) );
  or2 U2852 ( .A1(n2524), .A2(n1935), .Z(n2526) );
  inv1 U2853 ( .I(n2526), .ZN(n2602) );
  and2 U2854 ( .A1(n2525), .A2(n2602), .Z(n2528) );
  inv1 U2855 ( .I(n2525), .ZN(n2609) );
  and2 U2856 ( .A1(n2609), .A2(n2526), .Z(n2527) );
  or2 U2857 ( .A1(n2528), .A2(n2527), .Z(n460) );
  or2 U2859 ( .A1(n2529), .A2(n1937), .Z(n2530) );
  inv1 U2860 ( .I(n2530), .ZN(n2605) );
  and2 U2861 ( .A1(n463), .A2(n2605), .Z(n2533) );
  inv1 U2862 ( .I(n463), .ZN(n2531) );
  and2 U2863 ( .A1(n2531), .A2(n2530), .Z(n2532) );
  inv1 U2865 ( .I(n2534), .ZN(n3661) );
  and2 U2866 ( .A1(w4), .A2(f), .Z(n2536) );
  and2 U2867 ( .A1(g5), .A2(f), .Z(n2538) );
  and2 U2868 ( .A1(n), .A2(n2116), .Z(n2537) );
  or2 U2869 ( .A1(n2538), .A2(n2537), .Z(n2539) );
  and2 U2870 ( .A1(n2089), .A2(n2539), .Z(n2545) );
  inv1 U2871 ( .I(g5), .ZN(n2540) );
  and2 U2872 ( .A1(n2540), .A2(f), .Z(n2542) );
  and2 U2873 ( .A1(n439), .A2(n1928), .Z(n2541) );
  or2 U2874 ( .A1(n2542), .A2(n2541), .Z(n2543) );
  and2 U2875 ( .A1(n2581), .A2(n2543), .Z(n2544) );
  or2 U2876 ( .A1(n2545), .A2(n2544), .Z(n418) );
  and2 U2877 ( .A1(f5), .A2(f), .Z(n2546) );
  or2 U2878 ( .A1(n2546), .A2(n1949), .Z(n2548) );
  inv1 U2879 ( .I(n2548), .ZN(n2657) );
  and2 U2880 ( .A1(n2547), .A2(n2657), .Z(n2551) );
  and2 U2881 ( .A1(n2549), .A2(n2548), .Z(n2550) );
  or2 U2882 ( .A1(n2551), .A2(n2550), .Z(n417) );
  and2 U2883 ( .A1(n2552), .A2(n1920), .Z(n2555) );
  and2 U2884 ( .A1(n2553), .A2(n2058), .Z(n2554) );
  or2 U2885 ( .A1(n2555), .A2(n2554), .Z(n2558) );
  inv1 U2886 ( .I(n2558), .ZN(n2556) );
  and2 U2887 ( .A1(n2557), .A2(n2556), .Z(n2561) );
  and2 U2888 ( .A1(n2559), .A2(n2558), .Z(n2560) );
  or2 U2889 ( .A1(n2561), .A2(n2560), .Z(n414) );
  inv1 U2890 ( .I(n412), .ZN(n411) );
  and2 U2891 ( .A1(d5), .A2(f), .Z(n2562) );
  or2 U2892 ( .A1(n2562), .A2(n1929), .Z(n2564) );
  or2 U2894 ( .A1(n2563), .A2(n1927), .Z(n2565) );
  inv1 U2895 ( .I(n2565), .ZN(n2669) );
  and2 U2896 ( .A1(n2564), .A2(n2669), .Z(n2567) );
  inv1 U2897 ( .I(n2564), .ZN(n2660) );
  and2 U2898 ( .A1(n2660), .A2(n2565), .Z(n2566) );
  or2 U2899 ( .A1(n2567), .A2(n2566), .Z(n403) );
  and2 U2901 ( .A1(n406), .A2(n1913), .Z(n2573) );
  inv1 U2902 ( .I(n406), .ZN(n2571) );
  inv1 U2905 ( .I(n2574), .ZN(n3660) );
  or2 U2906 ( .A1(n2576), .A2(b6), .Z(n2575) );
  inv1 U2907 ( .I(n2575), .ZN(n3070) );
  and2 U2908 ( .A1(b6), .A2(n2576), .Z(n2577) );
  or2 U2909 ( .A1(n3070), .A2(n2577), .Z(n124) );
  or2 U2910 ( .A1(n2578), .A2(n3690), .Z(n3275) );
  inv1 U2911 ( .I(n3275), .ZN(n3277) );
  or2 U2912 ( .A1(n2579), .A2(z5), .Z(n3247) );
  inv1 U2913 ( .I(n3247), .ZN(n3249) );
  or2 U2914 ( .A1(n3277), .A2(n3249), .Z(n122) );
  inv1 U2915 ( .I(n122), .ZN(n3658) );
  inv1 U2916 ( .I(n124), .ZN(n3659) );
  inv1 U2917 ( .I(e6), .ZN(n2580) );
  or2 U2918 ( .A1(n2581), .A2(n2580), .Z(n2582) );
  or2 U2920 ( .A1(f), .A2(n2089), .Z(n2583) );
  or2 U2921 ( .A1(n2583), .A2(e6), .Z(n3592) );
  inv1 U2924 ( .I(x6), .ZN(n3643) );
  or2 U2925 ( .A1(n3579), .A2(n3643), .Z(n2936) );
  inv1 U2926 ( .I(n3579), .ZN(n2584) );
  or2 U2927 ( .A1(n2584), .A2(x6), .Z(n2585) );
  and2 U2928 ( .A1(n2936), .A2(n2585), .Z(d9) );
  and2 U2929 ( .A1(n1708), .A2(n3700), .Z(n3104) );
  or2 U2930 ( .A1(n3104), .A2(n3685), .Z(n3391) );
  inv1 U2931 ( .I(n3391), .ZN(n3393) );
  and2 U2932 ( .A1(n3684), .A2(n3393), .Z(n2714) );
  and2 U2933 ( .A1(p5), .A2(n2702), .Z(n2588) );
  and2 U2934 ( .A1(n3694), .A2(n2586), .Z(n2587) );
  or2 U2935 ( .A1(n2588), .A2(n2587), .Z(n3309) );
  or2 U2936 ( .A1(n2589), .A2(n3697), .Z(n3350) );
  or2 U2938 ( .A1(n2590), .A2(m5), .Z(n3324) );
  inv1 U2939 ( .I(n3324), .ZN(n3323) );
  and2 U2941 ( .A1(n5), .A2(n2703), .Z(n2593) );
  and2 U2942 ( .A1(n3696), .A2(n1992), .Z(n2592) );
  or2 U2943 ( .A1(n2593), .A2(n2592), .Z(n3306) );
  inv1 U2944 ( .I(n3306), .ZN(n3308) );
  and2 U2946 ( .A1(b1), .A2(n2594), .Z(n2596) );
  or2 U2949 ( .A1(n2596), .A2(n3048), .Z(n3313) );
  and2 U2950 ( .A1(o5), .A2(n2597), .Z(n2599) );
  or2 U2951 ( .A1(n2597), .A2(o5), .Z(n2598) );
  inv1 U2952 ( .I(n2598), .ZN(n3362) );
  or2 U2953 ( .A1(n2599), .A2(n3362), .Z(n3355) );
  or2 U2954 ( .A1(n3313), .A2(n3355), .Z(n2600) );
  or2 U2955 ( .A1(n3026), .A2(n2600), .Z(n2601) );
  inv1 U2956 ( .I(n2601), .ZN(n2695) );
  and2 U2957 ( .A1(r6), .A2(n2602), .Z(n2604) );
  or2 U2958 ( .A1(n2602), .A2(r6), .Z(n2603) );
  inv1 U2959 ( .I(n2603), .ZN(n3491) );
  and2 U2960 ( .A1(q6), .A2(n2605), .Z(n2607) );
  or2 U2961 ( .A1(n2605), .A2(q6), .Z(n2606) );
  inv1 U2962 ( .I(n2606), .ZN(n2614) );
  or2 U2963 ( .A1(n2608), .A2(o6), .Z(n3463) );
  and2 U2965 ( .A1(p6), .A2(n2609), .Z(n2611) );
  or2 U2966 ( .A1(n2609), .A2(p6), .Z(n2610) );
  inv1 U2967 ( .I(n2610), .ZN(n2612) );
  or2 U2971 ( .A1(n2615), .A2(n2614), .Z(n3483) );
  or2 U2972 ( .A1(n1920), .A2(n2617), .Z(n3548) );
  inv1 U2973 ( .I(n3548), .ZN(n3546) );
  or2 U2974 ( .A1(n2969), .A2(n3546), .Z(n3538) );
  inv1 U2978 ( .I(n2618), .ZN(n3098) );
  or2 U2979 ( .A1(n2026), .A2(n3098), .Z(n2620) );
  or2 U2981 ( .A1(n1909), .A2(n2621), .Z(n3505) );
  inv1 U2982 ( .I(n3505), .ZN(n3502) );
  or2 U2984 ( .A1(n3447), .A2(n3441), .Z(n3493) );
  or2 U2986 ( .A1(n3482), .A2(n3458), .Z(n3060) );
  and2 U2988 ( .A1(n2982), .A2(n1955), .Z(n2654) );
  and2 U2992 ( .A1(y5), .A2(n2651), .Z(n2629) );
  and2 U2993 ( .A1(n3691), .A2(n2627), .Z(n2628) );
  or2 U2994 ( .A1(n2629), .A2(n2628), .Z(n3189) );
  and2 U2996 ( .A1(x5), .A2(n2630), .Z(n2632) );
  or2 U2997 ( .A1(n2630), .A2(x5), .Z(n2631) );
  inv1 U2998 ( .I(n2631), .ZN(n3167) );
  or2 U2999 ( .A1(n3190), .A2(n3201), .Z(n2643) );
  or2 U3000 ( .A1(n2634), .A2(n2633), .Z(n3180) );
  or2 U3003 ( .A1(n1964), .A2(n2457), .Z(n2645) );
  inv1 U3004 ( .I(n2645), .ZN(n2639) );
  or2 U3005 ( .A1(n1965), .A2(v5), .Z(n2638) );
  inv1 U3006 ( .I(n2638), .ZN(n2646) );
  and2 U3009 ( .A1(w5), .A2(n2640), .Z(n2642) );
  or2 U3010 ( .A1(n2640), .A2(w5), .Z(n2641) );
  inv1 U3011 ( .I(n2641), .ZN(n2648) );
  or2 U3012 ( .A1(n3169), .A2(n3191), .Z(n3165) );
  or2 U3013 ( .A1(n2643), .A2(n3165), .Z(n3242) );
  or2 U3014 ( .A1(n2644), .A2(n3242), .Z(n3064) );
  and2 U3019 ( .A1(n2019), .A2(n3218), .Z(n2650) );
  or2 U3020 ( .A1(n2650), .A2(n3167), .Z(n3225) );
  and2 U3021 ( .A1(n3691), .A2(n2651), .Z(n2652) );
  or2 U3023 ( .A1(n2064), .A2(n2654), .Z(n2685) );
  or2 U3024 ( .A1(n2669), .A2(i6), .Z(n2655) );
  inv1 U3025 ( .I(n2655), .ZN(n2943) );
  and2 U3028 ( .A1(g6), .A2(n1913), .Z(n2656) );
  or2 U3029 ( .A1(n2056), .A2(n3643), .Z(n2918) );
  and2 U3030 ( .A1(f6), .A2(n2657), .Z(n2659) );
  or2 U3031 ( .A1(n2657), .A2(f6), .Z(n2658) );
  inv1 U3032 ( .I(n2658), .ZN(n2665) );
  and2 U3034 ( .A1(h6), .A2(n2660), .Z(n2661) );
  or2 U3037 ( .A1(n2662), .A2(n2918), .Z(n2663) );
  and2 U3038 ( .A1(n2664), .A2(n2663), .Z(n2668) );
  and2 U3044 ( .A1(i6), .A2(n2669), .Z(n2670) );
  and2 U3046 ( .A1(n2942), .A2(n2016), .Z(n2683) );
  and2 U3047 ( .A1(s6), .A2(n2673), .Z(n2674) );
  or2 U3048 ( .A1(n2673), .A2(s6), .Z(n2978) );
  and2 U3051 ( .A1(c6), .A2(n2675), .Z(n2677) );
  and2 U3052 ( .A1(n3687), .A2(n2687), .Z(n2676) );
  or2 U3053 ( .A1(n2677), .A2(n2676), .Z(n3259) );
  inv1 U3054 ( .I(n3259), .ZN(n3258) );
  or2 U3055 ( .A1(n3446), .A2(n3258), .Z(n2681) );
  or2 U3056 ( .A1(n124), .A2(n122), .Z(n3283) );
  and2 U3058 ( .A1(n3689), .A2(n2678), .Z(n2679) );
  or2 U3061 ( .A1(n3283), .A2(n3252), .Z(n3037) );
  or2 U3062 ( .A1(n2681), .A2(n3037), .Z(n2682) );
  or2 U3063 ( .A1(n2683), .A2(n2682), .Z(n2684) );
  or2 U3066 ( .A1(n2687), .A2(c6), .Z(n2688) );
  inv1 U3067 ( .I(n2688), .ZN(n3020) );
  and2 U3070 ( .A1(n3689), .A2(n2689), .Z(n2691) );
  or2 U3071 ( .A1(n3252), .A2(n3247), .Z(n3087) );
  inv1 U3072 ( .I(n3087), .ZN(n2690) );
  or2 U3073 ( .A1(n2691), .A2(n2690), .Z(n3248) );
  and2 U3077 ( .A1(n3256), .A2(n3037), .Z(n2693) );
  or2 U3078 ( .A1(n2693), .A2(n3258), .Z(n2993) );
  inv1 U3079 ( .I(n2993), .ZN(n2694) );
  and2 U3080 ( .A1(n2695), .A2(n2694), .Z(n2701) );
  and2 U3081 ( .A1(n2991), .A2(n3309), .Z(n2699) );
  or2 U3084 ( .A1(n3132), .A2(n2986), .Z(n3059) );
  or2 U3085 ( .A1(n2698), .A2(n3059), .Z(n2992) );
  and2 U3086 ( .A1(n2699), .A2(n2992), .Z(n2700) );
  and2 U3088 ( .A1(n3694), .A2(n2702), .Z(n2709) );
  inv1 U3089 ( .I(n3355), .ZN(n3361) );
  inv1 U3090 ( .I(n3313), .ZN(n3358) );
  and2 U3091 ( .A1(n3696), .A2(n2703), .Z(n2705) );
  or2 U3095 ( .A1(n2706), .A2(n3048), .Z(n3359) );
  and2 U3096 ( .A1(n3361), .A2(n3359), .Z(n2707) );
  or2 U3097 ( .A1(n2707), .A2(n3362), .Z(n3337) );
  and2 U3098 ( .A1(n3309), .A2(n3337), .Z(n2708) );
  or2 U3099 ( .A1(n2709), .A2(n2708), .Z(n2710) );
  and2 U3102 ( .A1(n2714), .A2(n3401), .Z(n2715) );
  or2 U3103 ( .A1(n2715), .A2(n3685), .Z(n2717) );
  or2 U3104 ( .A1(n2717), .A2(n2716), .Z(x9) );
  and2 U3105 ( .A1(n1052), .A2(n3698), .Z(n2718) );
  or2 U3106 ( .A1(n2718), .A2(n3700), .Z(n2719) );
  inv1 U3107 ( .I(n2719), .ZN(n2916) );
  and2 U3108 ( .A1(n1052), .A2(n3700), .Z(n2720) );
  inv1 U3109 ( .I(n2720), .ZN(n2724) );
  inv1 U3110 ( .I(n1355), .ZN(n2722) );
  inv1 U3111 ( .I(y6), .ZN(n2721) );
  or2 U3112 ( .A1(n2722), .A2(n2721), .Z(n2723) );
  and2 U3113 ( .A1(n2724), .A2(n2723), .Z(n2915) );
  or2 U3114 ( .A1(n2907), .A2(n840), .Z(n2912) );
  inv1 U3115 ( .I(n660), .ZN(n2725) );
  or2 U3116 ( .A1(n2726), .A2(n2725), .Z(n2886) );
  inv1 U3117 ( .I(n2886), .ZN(n2830) );
  inv1 U3118 ( .I(n1153), .ZN(n2728) );
  inv1 U3119 ( .I(n1148), .ZN(n2727) );
  or2 U3120 ( .A1(n2728), .A2(n2727), .Z(n2828) );
  and2 U3121 ( .A1(n2730), .A2(n2729), .Z(n2826) );
  or2 U3122 ( .A1(n2734), .A2(n2735), .Z(n2732) );
  and2 U3124 ( .A1(n2732), .A2(n2731), .Z(n2738) );
  inv1 U3125 ( .I(n683), .ZN(n2739) );
  inv1 U3126 ( .I(n2733), .ZN(n2740) );
  and2 U3127 ( .A1(n2739), .A2(n2740), .Z(n2737) );
  and2 U3128 ( .A1(n2735), .A2(n2734), .Z(n2736) );
  or2 U3129 ( .A1(n2737), .A2(n2736), .Z(n2819) );
  or2 U3130 ( .A1(n2738), .A2(n2819), .Z(n2742) );
  or2 U3131 ( .A1(n2740), .A2(n2739), .Z(n2741) );
  and2 U3132 ( .A1(n2742), .A2(n2741), .Z(n2744) );
  or2 U3133 ( .A1(n2745), .A2(n3671), .Z(n2743) );
  and2 U3134 ( .A1(n2744), .A2(n2743), .Z(n2748) );
  and2 U3135 ( .A1(n3672), .A2(n2749), .Z(n2747) );
  and2 U3136 ( .A1(n3671), .A2(n2745), .Z(n2746) );
  or2 U3137 ( .A1(n2747), .A2(n2746), .Z(n2818) );
  or2 U3138 ( .A1(n2748), .A2(n2818), .Z(n2751) );
  or2 U3139 ( .A1(n2749), .A2(n3672), .Z(n2750) );
  and2 U3140 ( .A1(n2751), .A2(n2750), .Z(n2824) );
  and2 U3141 ( .A1(n1930), .A2(n2793), .Z(n2752) );
  and2 U3142 ( .A1(n2792), .A2(n2752), .Z(n2755) );
  and2 U3143 ( .A1(n2790), .A2(n2791), .Z(n2754) );
  and2 U3144 ( .A1(n2786), .A2(n2787), .Z(n2753) );
  or2 U3145 ( .A1(n2754), .A2(n2753), .Z(n2797) );
  or2 U3146 ( .A1(n2755), .A2(n2797), .Z(n2760) );
  and2 U3147 ( .A1(n2761), .A2(n2762), .Z(n2757) );
  and2 U3148 ( .A1(n2784), .A2(n2785), .Z(n2756) );
  or2 U3149 ( .A1(n2757), .A2(n2756), .Z(n2801) );
  inv1 U3150 ( .I(w0), .ZN(n2758) );
  or2 U3151 ( .A1(n2801), .A2(n2758), .Z(n2759) );
  or2 U3152 ( .A1(n2760), .A2(n2759), .Z(n2764) );
  or2 U3153 ( .A1(n2762), .A2(n2761), .Z(n2763) );
  and2 U3154 ( .A1(n2764), .A2(n2763), .Z(n2805) );
  or2 U3155 ( .A1(n2766), .A2(n2765), .Z(n2767) );
  inv1 U3156 ( .I(n2767), .ZN(n2809) );
  or2 U3158 ( .A1(n2806), .A2(n2807), .Z(n2768) );
  and2 U3159 ( .A1(n2769), .A2(n2768), .Z(n2774) );
  and2 U3160 ( .A1(n2779), .A2(n2780), .Z(n2773) );
  or2 U3162 ( .A1(n2773), .A2(n2772), .Z(n2808) );
  or2 U3163 ( .A1(n2774), .A2(n2808), .Z(n2778) );
  or2 U3164 ( .A1(n2776), .A2(n2775), .Z(n2777) );
  and2 U3165 ( .A1(n2778), .A2(n2777), .Z(n2782) );
  or2 U3166 ( .A1(n2780), .A2(n2779), .Z(n2781) );
  and2 U3167 ( .A1(n2782), .A2(n2781), .Z(n2783) );
  or2 U3168 ( .A1(n2783), .A2(n2809), .Z(n2813) );
  or2 U3169 ( .A1(n2785), .A2(n2784), .Z(n2789) );
  or2 U3170 ( .A1(n2787), .A2(n2786), .Z(n2788) );
  and2 U3171 ( .A1(n2789), .A2(n2788), .Z(n2800) );
  or2 U3172 ( .A1(n2791), .A2(n2790), .Z(n2796) );
  or2 U3173 ( .A1(n2793), .A2(n2792), .Z(n2794) );
  or2 U3174 ( .A1(n2794), .A2(f), .Z(n2795) );
  and2 U3175 ( .A1(n2796), .A2(n2795), .Z(n2798) );
  or2 U3176 ( .A1(n2798), .A2(n2797), .Z(n2799) );
  and2 U3177 ( .A1(n2800), .A2(n2799), .Z(n2802) );
  or2 U3178 ( .A1(n2802), .A2(n2801), .Z(n2803) );
  and2 U3179 ( .A1(n2813), .A2(n2803), .Z(n2804) );
  and2 U3180 ( .A1(n2805), .A2(n2804), .Z(n2815) );
  and2 U3181 ( .A1(n2807), .A2(n2806), .Z(n2811) );
  or2 U3182 ( .A1(n2809), .A2(n2808), .Z(n2810) );
  or2 U3183 ( .A1(n2811), .A2(n2810), .Z(n2812) );
  and2 U3184 ( .A1(n2813), .A2(n2812), .Z(n2814) );
  or2 U3185 ( .A1(n2815), .A2(n2814), .Z(n2823) );
  and2 U3186 ( .A1(n2817), .A2(n2816), .Z(n2821) );
  or2 U3187 ( .A1(n2819), .A2(n2818), .Z(n2820) );
  or2 U3188 ( .A1(n2821), .A2(n2820), .Z(n2822) );
  or2 U3189 ( .A1(n2831), .A2(n2832), .Z(n2836) );
  inv1 U3190 ( .I(n2836), .ZN(n2825) );
  inv1 U3192 ( .I(n2829), .ZN(n2998) );
  and2 U3194 ( .A1(n2832), .A2(n2831), .Z(n2838) );
  and2 U3195 ( .A1(n719), .A2(n2833), .Z(n2834) );
  or2 U3196 ( .A1(n2834), .A2(n1146), .Z(n2835) );
  and2 U3197 ( .A1(n2836), .A2(n2835), .Z(n2837) );
  or2 U3198 ( .A1(n2838), .A2(n2837), .Z(n2997) );
  inv1 U3199 ( .I(n2997), .ZN(n2876) );
  or2 U3200 ( .A1(n2861), .A2(n3664), .Z(n2866) );
  or2 U3202 ( .A1(n2888), .A2(n2889), .Z(n2839) );
  or2 U3208 ( .A1(n2851), .A2(n3669), .Z(n2846) );
  and2 U3209 ( .A1(n2847), .A2(n2846), .Z(n2850) );
  or2 U3210 ( .A1(n2848), .A2(n3667), .Z(n2849) );
  and2 U3211 ( .A1(n2850), .A2(n2849), .Z(n2854) );
  and2 U3212 ( .A1(n3669), .A2(n2851), .Z(n2853) );
  and2 U3213 ( .A1(n3668), .A2(n2857), .Z(n2852) );
  or2 U3214 ( .A1(n2853), .A2(n2852), .Z(n2896) );
  or2 U3215 ( .A1(n2854), .A2(n2896), .Z(n2856) );
  or2 U3216 ( .A1(n2860), .A2(n3665), .Z(n2855) );
  or2 U3218 ( .A1(n2857), .A2(n3668), .Z(n2858) );
  and2 U3220 ( .A1(n3665), .A2(n2860), .Z(n2863) );
  and2 U3221 ( .A1(n3664), .A2(n2861), .Z(n2862) );
  or2 U3222 ( .A1(n2863), .A2(n2862), .Z(n2894) );
  or2 U3225 ( .A1(n2867), .A2(n666), .Z(n2868) );
  inv1 U3226 ( .I(n2868), .ZN(n2891) );
  or2 U3228 ( .A1(n2870), .A2(n3666), .Z(n2871) );
  and2 U3229 ( .A1(n2872), .A2(n2871), .Z(n2875) );
  or2 U3230 ( .A1(n2873), .A2(n660), .Z(n2874) );
  inv1 U3231 ( .I(n2874), .ZN(n2890) );
  and2 U3233 ( .A1(n2876), .A2(n2887), .Z(n2877) );
  or2 U3237 ( .A1(n2101), .A2(n812), .Z(n2882) );
  and2 U3238 ( .A1(n2883), .A2(n2882), .Z(n2884) );
  and2 U3240 ( .A1(n1063), .A2(n1067), .Z(n2904) );
  and2 U3242 ( .A1(n2889), .A2(n2888), .Z(n2893) );
  or2 U3243 ( .A1(n2891), .A2(n2890), .Z(n2892) );
  or2 U3244 ( .A1(n2893), .A2(n2892), .Z(n2899) );
  or2 U3245 ( .A1(n2895), .A2(n2894), .Z(n2897) );
  or2 U3246 ( .A1(n2897), .A2(n2896), .Z(n2898) );
  or2 U3247 ( .A1(n2899), .A2(n2898), .Z(n2900) );
  inv1 U3249 ( .I(n2902), .ZN(n2903) );
  and2 U3251 ( .A1(n840), .A2(n2907), .Z(n2910) );
  and2 U3252 ( .A1(n841), .A2(n2908), .Z(n2909) );
  or2 U3253 ( .A1(n2910), .A2(n2909), .Z(n2911) );
  or2 U3254 ( .A1(n2911), .A2(n1061), .Z(n2913) );
  and2 U3255 ( .A1(n2913), .A2(n2912), .Z(n2914) );
  inv1 U3257 ( .I(n2918), .ZN(n2919) );
  and2 U3258 ( .A1(n3625), .A2(n2919), .Z(n2920) );
  or2 U3259 ( .A1(n2920), .A2(n2002), .Z(n2927) );
  inv1 U3260 ( .I(n2927), .ZN(n2921) );
  or2 U3261 ( .A1(n2921), .A2(n1923), .Z(n2929) );
  inv1 U3262 ( .I(n2929), .ZN(n2922) );
  or2 U3263 ( .A1(n2922), .A2(n3617), .Z(n2923) );
  or2 U3264 ( .A1(n2923), .A2(n1981), .Z(n2926) );
  inv1 U3265 ( .I(n2923), .ZN(n2924) );
  or2 U3266 ( .A1(n2924), .A2(n3575), .Z(n2925) );
  and2 U3267 ( .A1(n2926), .A2(n2925), .Z(i9) );
  inv1 U3268 ( .I(n1923), .ZN(n3616) );
  or2 U3269 ( .A1(n2927), .A2(n3616), .Z(n2928) );
  and2 U3270 ( .A1(n2929), .A2(n2928), .Z(j9) );
  inv1 U3271 ( .I(n3626), .ZN(n3595) );
  and2 U3272 ( .A1(n2057), .A2(n3595), .Z(n2931) );
  or2 U3273 ( .A1(n3578), .A2(n2936), .Z(n2930) );
  and2 U3274 ( .A1(n2931), .A2(n2930), .Z(n2935) );
  and2 U3275 ( .A1(x6), .A2(n3625), .Z(n2932) );
  or2 U3276 ( .A1(n2932), .A2(n3626), .Z(n2933) );
  and2 U3277 ( .A1(n2056), .A2(n2933), .Z(n2934) );
  or2 U3278 ( .A1(n2935), .A2(n2934), .Z(k9) );
  inv1 U3279 ( .I(n2936), .ZN(n2937) );
  or2 U3280 ( .A1(n2937), .A2(n3591), .Z(n2938) );
  or2 U3281 ( .A1(n2938), .A2(n2070), .Z(n2941) );
  inv1 U3282 ( .I(n2938), .ZN(n2939) );
  or2 U3283 ( .A1(n2939), .A2(n3578), .Z(n2940) );
  and2 U3284 ( .A1(n2941), .A2(n2940), .Z(l9) );
  inv1 U3285 ( .I(n3647), .ZN(n3649) );
  and2 U3286 ( .A1(n2944), .A2(n3649), .Z(n2956) );
  inv1 U3287 ( .I(n2945), .ZN(n2946) );
  or2 U3288 ( .A1(n2946), .A2(n2957), .Z(n3561) );
  inv1 U3289 ( .I(n3561), .ZN(n3563) );
  or2 U3290 ( .A1(n3563), .A2(n1919), .Z(n2963) );
  inv1 U3291 ( .I(n2963), .ZN(n2948) );
  or2 U3292 ( .A1(n2948), .A2(n2947), .Z(n2951) );
  or2 U3293 ( .A1(n2951), .A2(n2949), .Z(n2950) );
  and2 U3294 ( .A1(n3647), .A2(n2950), .Z(n2954) );
  inv1 U3295 ( .I(n2951), .ZN(n2952) );
  or2 U3296 ( .A1(n2952), .A2(n3554), .Z(n2953) );
  and2 U3297 ( .A1(n2954), .A2(n2953), .Z(n2955) );
  or2 U3298 ( .A1(n2956), .A2(n2955), .Z(m9) );
  inv1 U3299 ( .I(n1919), .ZN(n3532) );
  or2 U3300 ( .A1(n2957), .A2(n3532), .Z(n2958) );
  and2 U3301 ( .A1(n3649), .A2(n2958), .Z(n2959) );
  and2 U3302 ( .A1(n2960), .A2(n2959), .Z(n2965) );
  or2 U3303 ( .A1(n3561), .A2(n3532), .Z(n2961) );
  and2 U3304 ( .A1(n3647), .A2(n2961), .Z(n2962) );
  and2 U3305 ( .A1(n2963), .A2(n2962), .Z(n2964) );
  or2 U3306 ( .A1(n2965), .A2(n2964), .Z(n9) );
  or2 U3307 ( .A1(n2028), .A2(n3548), .Z(n2966) );
  and2 U3308 ( .A1(n3647), .A2(n2966), .Z(n2968) );
  or2 U3309 ( .A1(n3531), .A2(n3546), .Z(n2967) );
  and2 U3310 ( .A1(n2968), .A2(n2967), .Z(n2975) );
  and2 U3311 ( .A1(n2969), .A2(n3531), .Z(n2972) );
  and2 U3312 ( .A1(n2970), .A2(n2028), .Z(n2971) );
  or2 U3313 ( .A1(n2972), .A2(n2971), .Z(n2973) );
  and2 U3314 ( .A1(n3649), .A2(n2973), .Z(n2974) );
  or2 U3315 ( .A1(n2975), .A2(n2974), .Z(o9) );
  inv1 U3316 ( .I(n3538), .ZN(n3535) );
  or2 U3317 ( .A1(n3647), .A2(n3535), .Z(n2977) );
  or2 U3318 ( .A1(n3649), .A2(n3538), .Z(n2976) );
  and2 U3319 ( .A1(n2977), .A2(n2976), .Z(p9) );
  and2 U3320 ( .A1(n2978), .A2(n3446), .Z(n2980) );
  or2 U3321 ( .A1(n2980), .A2(n2979), .Z(n2981) );
  inv1 U3322 ( .I(n2981), .ZN(n2985) );
  or2 U3326 ( .A1(n2061), .A2(n3183), .Z(n3013) );
  or2 U3328 ( .A1(n2059), .A2(n3185), .Z(n2990) );
  and2 U3329 ( .A1(n3013), .A2(n2990), .Z(u9) );
  inv1 U3336 ( .I(n3314), .ZN(n3312) );
  or2 U3337 ( .A1(n3407), .A2(n3312), .Z(n2996) );
  and2 U3338 ( .A1(n3053), .A2(n2996), .Z(v9) );
  or2 U3339 ( .A1(n2998), .A2(n2997), .Z(w9) );
  or2 U3340 ( .A1(n2061), .A2(n3169), .Z(n2999) );
  inv1 U3345 ( .I(n3002), .ZN(n3001) );
  and2 U3347 ( .A1(n3002), .A2(n3190), .Z(n3003) );
  or2 U3348 ( .A1(n3004), .A2(n3003), .Z(y9) );
  or2 U3349 ( .A1(n3005), .A2(n2019), .Z(n3006) );
  and2 U3350 ( .A1(n3007), .A2(n3006), .Z(z9) );
  or2 U3351 ( .A1(n3008), .A2(n3217), .Z(n3009) );
  or2 U3352 ( .A1(n3009), .A2(n2068), .Z(n3012) );
  inv1 U3353 ( .I(n3009), .ZN(n3010) );
  or2 U3354 ( .A1(n3010), .A2(n3191), .Z(n3011) );
  and2 U3355 ( .A1(n3012), .A2(n3011), .Z(a10) );
  inv1 U3356 ( .I(n3013), .ZN(n3014) );
  or2 U3357 ( .A1(n3014), .A2(n2014), .Z(n3015) );
  inv1 U3358 ( .I(n3186), .ZN(n3184) );
  or2 U3359 ( .A1(n3015), .A2(n3184), .Z(n3018) );
  inv1 U3360 ( .I(n3015), .ZN(n3016) );
  or2 U3361 ( .A1(n3016), .A2(n3186), .Z(n3017) );
  and2 U3362 ( .A1(n3018), .A2(n3017), .Z(b10) );
  or2 U3363 ( .A1(n3048), .A2(n3358), .Z(n3019) );
  and2 U3364 ( .A1(n3361), .A2(n3019), .Z(n3031) );
  or2 U3365 ( .A1(n3370), .A2(n3020), .Z(n3021) );
  or2 U3366 ( .A1(n3048), .A2(n3021), .Z(n3025) );
  or2 U3368 ( .A1(n3025), .A2(n3024), .Z(n3029) );
  or2 U3370 ( .A1(n3048), .A2(n3370), .Z(n3027) );
  or2 U3371 ( .A1(n3371), .A2(n3027), .Z(n3028) );
  and2 U3372 ( .A1(n3029), .A2(n3028), .Z(n3030) );
  inv1 U3375 ( .I(n3034), .ZN(n3033) );
  and2 U3376 ( .A1(n3309), .A2(n3033), .Z(n3036) );
  inv1 U3377 ( .I(n3309), .ZN(n3307) );
  and2 U3378 ( .A1(n3307), .A2(n3034), .Z(n3035) );
  inv1 U3380 ( .I(n3037), .ZN(n3038) );
  or2 U3382 ( .A1(n3059), .A2(n3079), .Z(n3039) );
  and2 U3385 ( .A1(n3259), .A2(n3042), .Z(n3043) );
  and2 U3386 ( .A1(n3371), .A2(n3043), .Z(n3047) );
  and2 U3390 ( .A1(n3049), .A2(n3050), .Z(d10) );
  or2 U3391 ( .A1(n3051), .A2(n3358), .Z(n3052) );
  and2 U3392 ( .A1(n1917), .A2(n3052), .Z(e10) );
  inv1 U3393 ( .I(n3053), .ZN(n3054) );
  or2 U3394 ( .A1(n3054), .A2(n3323), .Z(n3056) );
  or2 U3395 ( .A1(n3056), .A2(n3308), .Z(n3055) );
  inv1 U3396 ( .I(n3055), .ZN(n3058) );
  and2 U3397 ( .A1(n3308), .A2(n3056), .Z(n3057) );
  or2 U3398 ( .A1(n3058), .A2(n3057), .Z(f10) );
  inv1 U3399 ( .I(n3059), .ZN(n3063) );
  or2 U3400 ( .A1(n3060), .A2(n2041), .Z(n3061) );
  and2 U3401 ( .A1(n3063), .A2(n3131), .Z(n3065) );
  and2 U3403 ( .A1(n3258), .A2(n3253), .Z(n3067) );
  and2 U3404 ( .A1(n3259), .A2(n3256), .Z(n3066) );
  or2 U3405 ( .A1(n3067), .A2(n3066), .Z(n3068) );
  and2 U3406 ( .A1(n2062), .A2(n3068), .Z(n3078) );
  and2 U3407 ( .A1(n3658), .A2(n3255), .Z(n3069) );
  or2 U3408 ( .A1(n3069), .A2(n3248), .Z(n3276) );
  and2 U3409 ( .A1(n3659), .A2(n3276), .Z(n3071) );
  or2 U3410 ( .A1(n3071), .A2(n3070), .Z(n3072) );
  and2 U3411 ( .A1(n3258), .A2(n3072), .Z(n3075) );
  inv1 U3412 ( .I(n3072), .ZN(n3073) );
  and2 U3413 ( .A1(n3259), .A2(n3073), .Z(n3074) );
  or2 U3414 ( .A1(n3075), .A2(n3074), .Z(n3076) );
  and2 U3415 ( .A1(n3095), .A2(n3076), .Z(n3077) );
  or2 U3416 ( .A1(n3078), .A2(n3077), .Z(i10) );
  inv1 U3417 ( .I(n3248), .ZN(n3246) );
  inv1 U3418 ( .I(n3079), .ZN(n3243) );
  and2 U3419 ( .A1(n3246), .A2(n3243), .Z(n3080) );
  inv1 U3421 ( .I(n3276), .ZN(n3274) );
  inv1 U3425 ( .I(n3084), .ZN(n3085) );
  or2 U3426 ( .A1(n3086), .A2(n3085), .Z(j10) );
  or2 U3428 ( .A1(n3255), .A2(n3249), .Z(n3088) );
  and2 U3430 ( .A1(n3275), .A2(n3252), .Z(n3091) );
  and2 U3431 ( .A1(n3277), .A2(n3255), .Z(n3090) );
  or2 U3432 ( .A1(n3091), .A2(n3090), .Z(n3092) );
  and2 U3433 ( .A1(n3095), .A2(n3092), .Z(n3093) );
  or2 U3434 ( .A1(n3094), .A2(n3093), .Z(k10) );
  or2 U3435 ( .A1(n3095), .A2(n3658), .Z(n3097) );
  or2 U3436 ( .A1(n2062), .A2(n122), .Z(n3096) );
  and2 U3437 ( .A1(n3097), .A2(n3096), .Z(l10) );
  or2 U3439 ( .A1(n2060), .A2(n3447), .Z(n3125) );
  inv1 U3440 ( .I(n3447), .ZN(n3445) );
  or2 U3441 ( .A1(n2042), .A2(n3445), .Z(n3100) );
  and2 U3442 ( .A1(n3125), .A2(n3100), .Z(m10) );
  and2 U3444 ( .A1(n3684), .A2(n3705), .Z(n3102) );
  and2 U3445 ( .A1(n19), .A2(n3685), .Z(n3101) );
  or2 U3446 ( .A1(n3102), .A2(n3101), .Z(n3103) );
  and2 U3447 ( .A1(n3403), .A2(n3103), .Z(n3109) );
  and2 U3448 ( .A1(n19), .A2(n3104), .Z(n3107) );
  inv1 U3449 ( .I(n3104), .ZN(n3105) );
  and2 U3450 ( .A1(n3684), .A2(n3105), .Z(n3106) );
  or2 U3451 ( .A1(n3107), .A2(n3106), .Z(n3392) );
  inv1 U3452 ( .I(n3392), .ZN(n3390) );
  and2 U3453 ( .A1(n3401), .A2(n3390), .Z(n3108) );
  or2 U3454 ( .A1(n3109), .A2(n3108), .Z(z850) );
  and2 U3455 ( .A1(n3393), .A2(n3401), .Z(n3111) );
  and2 U3456 ( .A1(n3391), .A2(n3403), .Z(n3110) );
  or2 U3457 ( .A1(n3111), .A2(n3110), .Z(n3112) );
  inv1 U3458 ( .I(n3112), .ZN(p10) );
  and2 U3461 ( .A1(n1988), .A2(n3120), .Z(n3114) );
  or2 U3462 ( .A1(n3114), .A2(n2008), .Z(n3117) );
  or2 U3464 ( .A1(n2038), .A2(n3448), .Z(n3116) );
  and2 U3466 ( .A1(n3116), .A2(n3115), .Z(r10) );
  or2 U3467 ( .A1(n3117), .A2(n1995), .Z(n3118) );
  and2 U3468 ( .A1(n3119), .A2(n3118), .Z(s10) );
  or2 U3469 ( .A1(n3120), .A2(n2074), .Z(n3121) );
  or2 U3470 ( .A1(n3121), .A2(n1988), .Z(n3124) );
  inv1 U3471 ( .I(n3121), .ZN(n3122) );
  or2 U3472 ( .A1(n3122), .A2(n3442), .Z(n3123) );
  and2 U3473 ( .A1(n3124), .A2(n3123), .Z(t10) );
  inv1 U3474 ( .I(n3125), .ZN(n3126) );
  or2 U3475 ( .A1(n3126), .A2(n3462), .Z(n3127) );
  or2 U3476 ( .A1(n3127), .A2(n2021), .Z(n3130) );
  inv1 U3477 ( .I(n3127), .ZN(n3128) );
  or2 U3478 ( .A1(n3128), .A2(n3441), .Z(n3129) );
  and2 U3479 ( .A1(n3130), .A2(n3129), .Z(u10) );
  and2 U3480 ( .A1(n3683), .A2(n2024), .Z(n3144) );
  and2 U3481 ( .A1(n3418), .A2(n3133), .Z(n3135) );
  or2 U3482 ( .A1(n3135), .A2(n3134), .Z(n3138) );
  or2 U3483 ( .A1(n3138), .A2(n3136), .Z(n3137) );
  and2 U3484 ( .A1(n3522), .A2(n3137), .Z(n3142) );
  inv1 U3485 ( .I(n3138), .ZN(n3140) );
  or2 U3486 ( .A1(n3140), .A2(n3139), .Z(n3141) );
  and2 U3487 ( .A1(n3142), .A2(n3141), .Z(n3143) );
  or2 U3488 ( .A1(n3144), .A2(n3143), .Z(v10) );
  and2 U3489 ( .A1(n3145), .A2(n2024), .Z(n3147) );
  or2 U3490 ( .A1(n3147), .A2(n3146), .Z(n3149) );
  inv1 U3491 ( .I(n3149), .ZN(n3148) );
  and2 U3493 ( .A1(n3418), .A2(n3149), .Z(n3150) );
  or2 U3494 ( .A1(n3151), .A2(n3150), .Z(w10) );
  and2 U3495 ( .A1(n3152), .A2(n3423), .Z(n3154) );
  and2 U3496 ( .A1(n1983), .A2(n3426), .Z(n3153) );
  or2 U3497 ( .A1(n3154), .A2(n3153), .Z(n3155) );
  and2 U3498 ( .A1(n2024), .A2(n3155), .Z(n3162) );
  or2 U3499 ( .A1(n3423), .A2(n3156), .Z(n3157) );
  and2 U3500 ( .A1(n3522), .A2(n3157), .Z(n3160) );
  or2 U3501 ( .A1(n3426), .A2(n3158), .Z(n3159) );
  and2 U3502 ( .A1(n3160), .A2(n3159), .Z(n3161) );
  or2 U3503 ( .A1(n3162), .A2(n3161), .Z(x10) );
  or2 U3504 ( .A1(n3522), .A2(n3419), .Z(n3164) );
  or2 U3505 ( .A1(n2024), .A2(n3417), .Z(n3163) );
  and2 U3506 ( .A1(n3164), .A2(n3163), .Z(y10) );
  inv1 U3507 ( .I(n3165), .ZN(n3166) );
  and2 U3509 ( .A1(n2019), .A2(n3206), .Z(n3168) );
  or2 U3510 ( .A1(n3168), .A2(n3167), .Z(n3172) );
  inv1 U3511 ( .I(n3169), .ZN(n3170) );
  or2 U3512 ( .A1(n3170), .A2(n3217), .Z(n3173) );
  inv1 U3513 ( .I(n3173), .ZN(n3171) );
  and2 U3516 ( .A1(n3174), .A2(n3173), .Z(n3175) );
  and2 U3518 ( .A1(n3177), .A2(n3178), .Z(n3182) );
  or2 U3521 ( .A1(n3182), .A2(n3181), .Z(n3213) );
  inv1 U3522 ( .I(n3213), .ZN(n3209) );
  and2 U3524 ( .A1(n3186), .A2(n3185), .Z(n3187) );
  or2 U3525 ( .A1(n3188), .A2(n3187), .Z(n3195) );
  and2 U3526 ( .A1(n2068), .A2(n3189), .Z(n3193) );
  or2 U3528 ( .A1(n3193), .A2(n3192), .Z(n3196) );
  inv1 U3529 ( .I(n3196), .ZN(n3194) );
  and2 U3530 ( .A1(n3195), .A2(n3194), .Z(n3199) );
  inv1 U3531 ( .I(n3195), .ZN(n3197) );
  and2 U3532 ( .A1(n3197), .A2(n3196), .Z(n3198) );
  inv1 U3534 ( .I(n3202), .ZN(n3200) );
  and2 U3535 ( .A1(n3201), .A2(n3200), .Z(n3204) );
  and2 U3536 ( .A1(n2019), .A2(n3202), .Z(n3203) );
  inv1 U3538 ( .I(n1963), .ZN(n3205) );
  and2 U3539 ( .A1(n3228), .A2(n3205), .Z(n3208) );
  and2 U3541 ( .A1(n3229), .A2(n1963), .Z(n3207) );
  or2 U3542 ( .A1(n3208), .A2(n3207), .Z(n3212) );
  inv1 U3546 ( .I(n3225), .ZN(n3222) );
  inv1 U3547 ( .I(n3218), .ZN(n3216) );
  and2 U3548 ( .A1(n3217), .A2(n3216), .Z(n3221) );
  inv1 U3549 ( .I(n3217), .ZN(n3219) );
  and2 U3550 ( .A1(n3219), .A2(n3218), .Z(n3220) );
  or2 U3551 ( .A1(n3221), .A2(n3220), .Z(n3223) );
  and2 U3552 ( .A1(n3222), .A2(n3223), .Z(n3227) );
  inv1 U3553 ( .I(n3223), .ZN(n3224) );
  and2 U3554 ( .A1(n3225), .A2(n3224), .Z(n3226) );
  or2 U3555 ( .A1(n3227), .A2(n3226), .Z(n3237) );
  inv1 U3556 ( .I(n3237), .ZN(n3233) );
  and2 U3557 ( .A1(n2014), .A2(n3228), .Z(n3232) );
  inv1 U3562 ( .I(n3235), .ZN(n3236) );
  or2 U3563 ( .A1(n3237), .A2(n3236), .Z(n3238) );
  and2 U3564 ( .A1(n3239), .A2(n3238), .Z(n3240) );
  and2 U3567 ( .A1(n3243), .A2(n3242), .Z(n3245) );
  and2 U3568 ( .A1(n2061), .A2(n3243), .Z(n3244) );
  or2 U3569 ( .A1(n3245), .A2(n3244), .Z(n3273) );
  and2 U3570 ( .A1(n3247), .A2(n3246), .Z(n3251) );
  and2 U3571 ( .A1(n3249), .A2(n3248), .Z(n3250) );
  or2 U3572 ( .A1(n3251), .A2(n3250), .Z(n3270) );
  inv1 U3573 ( .I(n3270), .ZN(n3266) );
  or2 U3574 ( .A1(n3253), .A2(n3252), .Z(n3254) );
  inv1 U3575 ( .I(n3254), .ZN(n3282) );
  or2 U3576 ( .A1(n3256), .A2(n3255), .Z(n3257) );
  inv1 U3577 ( .I(n3257), .ZN(n3284) );
  or2 U3578 ( .A1(n3282), .A2(n3284), .Z(n3263) );
  inv1 U3579 ( .I(n3263), .ZN(n3280) );
  and2 U3580 ( .A1(n118), .A2(n3258), .Z(n3262) );
  inv1 U3581 ( .I(n118), .ZN(n3260) );
  and2 U3582 ( .A1(n3260), .A2(n3259), .Z(n3261) );
  or2 U3583 ( .A1(n3262), .A2(n3261), .Z(n3295) );
  and2 U3584 ( .A1(n3280), .A2(n3295), .Z(n3265) );
  inv1 U3585 ( .I(n3295), .ZN(n3290) );
  and2 U3586 ( .A1(n3263), .A2(n3290), .Z(n3264) );
  or2 U3587 ( .A1(n3265), .A2(n3264), .Z(n3268) );
  inv1 U3590 ( .I(n3268), .ZN(n3269) );
  or2 U3591 ( .A1(n3270), .A2(n3269), .Z(n3271) );
  and2 U3594 ( .A1(n3275), .A2(n3274), .Z(n3279) );
  and2 U3595 ( .A1(n3277), .A2(n3276), .Z(n3278) );
  or2 U3596 ( .A1(n3279), .A2(n3278), .Z(n3281) );
  and2 U3597 ( .A1(n3281), .A2(n3280), .Z(n3289) );
  inv1 U3598 ( .I(n3281), .ZN(n3287) );
  and2 U3599 ( .A1(n3283), .A2(n3282), .Z(n3285) );
  or2 U3600 ( .A1(n3285), .A2(n3284), .Z(n3286) );
  inv1 U3605 ( .I(n3293), .ZN(n3294) );
  or2 U3606 ( .A1(n3295), .A2(n3294), .Z(n3296) );
  or2 U3609 ( .A1(n3301), .A2(n3300), .Z(n3305) );
  or2 U3611 ( .A1(n3303), .A2(n3302), .Z(n3304) );
  and2 U3613 ( .A1(n3307), .A2(n3306), .Z(n3311) );
  and2 U3614 ( .A1(n3309), .A2(n3308), .Z(n3310) );
  or2 U3615 ( .A1(n3311), .A2(n3310), .Z(n3318) );
  and2 U3616 ( .A1(n3313), .A2(n3312), .Z(n3316) );
  or2 U3618 ( .A1(n3316), .A2(n3315), .Z(n3319) );
  inv1 U3619 ( .I(n3319), .ZN(n3317) );
  inv1 U3621 ( .I(n3318), .ZN(n3320) );
  and2 U3624 ( .A1(n3323), .A2(n3347), .Z(n3326) );
  inv1 U3625 ( .I(n3347), .ZN(n3349) );
  and2 U3628 ( .A1(n3361), .A2(n3327), .Z(n3330) );
  inv1 U3629 ( .I(n3327), .ZN(n3328) );
  and2 U3630 ( .A1(n3355), .A2(n3328), .Z(n3329) );
  or2 U3631 ( .A1(n3330), .A2(n3329), .Z(n3341) );
  inv1 U3632 ( .I(n3337), .ZN(n3334) );
  inv1 U3633 ( .I(n3359), .ZN(n3331) );
  and2 U3634 ( .A1(n3370), .A2(n3331), .Z(n3333) );
  and2 U3635 ( .A1(n1997), .A2(n3359), .Z(n3332) );
  or2 U3636 ( .A1(n3333), .A2(n3332), .Z(n3335) );
  and2 U3637 ( .A1(n3334), .A2(n3335), .Z(n3339) );
  inv1 U3638 ( .I(n3335), .ZN(n3336) );
  and2 U3639 ( .A1(n3337), .A2(n3336), .Z(n3338) );
  or2 U3640 ( .A1(n3339), .A2(n3338), .Z(n3342) );
  inv1 U3641 ( .I(n3342), .ZN(n3340) );
  inv1 U3646 ( .I(n3408), .ZN(n3346) );
  and2 U3648 ( .A1(n3348), .A2(n3347), .Z(n3352) );
  and2 U3649 ( .A1(n3350), .A2(n3349), .Z(n3351) );
  or2 U3650 ( .A1(n3352), .A2(n3351), .Z(n3353) );
  and2 U3651 ( .A1(n3361), .A2(n3353), .Z(n3357) );
  inv1 U3652 ( .I(n3353), .ZN(n3354) );
  inv1 U3658 ( .I(n3366), .ZN(n3364) );
  and2 U3659 ( .A1(n1991), .A2(n3364), .Z(n3369) );
  inv1 U3660 ( .I(n1991), .ZN(n3367) );
  and2 U3661 ( .A1(n3367), .A2(n3366), .Z(n3368) );
  or2 U3663 ( .A1(n3371), .A2(n3370), .Z(n3374) );
  inv1 U3664 ( .I(n3374), .ZN(n3372) );
  inv1 U3671 ( .I(n3379), .ZN(n3381) );
  inv1 U3674 ( .I(n3410), .ZN(n3384) );
  and2 U3677 ( .A1(n1701), .A2(n3393), .Z(n3389) );
  inv1 U3678 ( .I(n1701), .ZN(n3387) );
  and2 U3679 ( .A1(n3387), .A2(n3391), .Z(n3388) );
  or2 U3680 ( .A1(n3389), .A2(n3388), .Z(n3400) );
  and2 U3682 ( .A1(n3391), .A2(n3390), .Z(n3395) );
  and2 U3683 ( .A1(n3393), .A2(n3392), .Z(n3394) );
  or2 U3684 ( .A1(n3395), .A2(n3394), .Z(n3404) );
  and2 U3685 ( .A1(n3397), .A2(n3396), .Z(n3398) );
  inv1 U3687 ( .I(n3400), .ZN(n3402) );
  or2 U3688 ( .A1(n3401), .A2(n3402), .Z(n3406) );
  or2 U3694 ( .A1(n3414), .A2(n3413), .Z(n3415) );
  and2 U3695 ( .A1(n3416), .A2(n3415), .Z(a11) );
  and2 U3696 ( .A1(n3418), .A2(n3417), .Z(n3422) );
  and2 U3697 ( .A1(n3420), .A2(n3419), .Z(n3421) );
  or2 U3698 ( .A1(n3422), .A2(n3421), .Z(n3424) );
  and2 U3699 ( .A1(n3423), .A2(n3424), .Z(n3428) );
  inv1 U3700 ( .I(n3424), .ZN(n3425) );
  and2 U3701 ( .A1(n3426), .A2(n3425), .Z(n3427) );
  or2 U3702 ( .A1(n3428), .A2(n3427), .Z(n3434) );
  inv1 U3703 ( .I(n3434), .ZN(n3433) );
  and2 U3704 ( .A1(n1584), .A2(n3433), .Z(n3431) );
  inv1 U3705 ( .I(n1584), .ZN(n3429) );
  and2 U3706 ( .A1(n3429), .A2(n3434), .Z(n3430) );
  or2 U3707 ( .A1(n3431), .A2(n3430), .Z(n3523) );
  inv1 U3708 ( .I(n3523), .ZN(n3432) );
  or2 U3709 ( .A1(n3432), .A2(n3522), .Z(n3440) );
  and2 U3710 ( .A1(n1564), .A2(n3433), .Z(n3437) );
  inv1 U3711 ( .I(n1564), .ZN(n3435) );
  and2 U3712 ( .A1(n3435), .A2(n3434), .Z(n3436) );
  or2 U3713 ( .A1(n3437), .A2(n3436), .Z(n3524) );
  inv1 U3714 ( .I(n3524), .ZN(n3438) );
  or2 U3715 ( .A1(n3438), .A2(n2024), .Z(n3439) );
  and2 U3716 ( .A1(n3440), .A2(n3439), .Z(n3517) );
  and2 U3718 ( .A1(n3442), .A2(n2021), .Z(n3443) );
  or2 U3719 ( .A1(n3444), .A2(n3443), .Z(n3452) );
  and2 U3721 ( .A1(n3448), .A2(n3447), .Z(n3449) );
  or2 U3722 ( .A1(n3450), .A2(n3449), .Z(n3453) );
  inv1 U3723 ( .I(n3453), .ZN(n3451) );
  and2 U3724 ( .A1(n3452), .A2(n3451), .Z(n3456) );
  inv1 U3725 ( .I(n3452), .ZN(n3454) );
  and2 U3726 ( .A1(n3454), .A2(n3453), .Z(n3455) );
  inv1 U3728 ( .I(n3459), .ZN(n3457) );
  and2 U3729 ( .A1(n3458), .A2(n3457), .Z(n3461) );
  and2 U3730 ( .A1(n1995), .A2(n3459), .Z(n3460) );
  inv1 U3736 ( .I(n3483), .ZN(n3466) );
  and2 U3737 ( .A1(n2074), .A2(n3466), .Z(n3469) );
  inv1 U3738 ( .I(n3494), .ZN(n3467) );
  and2 U3739 ( .A1(n3467), .A2(n2008), .Z(n3468) );
  or2 U3740 ( .A1(n3469), .A2(n3468), .Z(n3470) );
  and2 U3741 ( .A1(n1955), .A2(n3470), .Z(n3474) );
  inv1 U3742 ( .I(n3470), .ZN(n3471) );
  and2 U3743 ( .A1(n2078), .A2(n3471), .Z(n3473) );
  or2 U3744 ( .A1(n3474), .A2(n3473), .Z(n3477) );
  inv1 U3745 ( .I(n3477), .ZN(n3475) );
  and2 U3746 ( .A1(n3476), .A2(n3475), .Z(n3480) );
  inv1 U3747 ( .I(n3476), .ZN(n3478) );
  or2 U3751 ( .A1(n3481), .A2(n2042), .Z(n3515) );
  inv1 U3752 ( .I(n3482), .ZN(n3484) );
  or2 U3753 ( .A1(n3484), .A2(n3483), .Z(n3490) );
  inv1 U3754 ( .I(n2007), .ZN(n3485) );
  or2 U3757 ( .A1(n3489), .A2(n3488), .Z(n3509) );
  and2 U3758 ( .A1(n3490), .A2(n1995), .Z(n3492) );
  or2 U3759 ( .A1(n3492), .A2(n3491), .Z(n3497) );
  inv1 U3760 ( .I(n3493), .ZN(n3495) );
  or2 U3761 ( .A1(n3495), .A2(n2074), .Z(n3498) );
  inv1 U3762 ( .I(n3498), .ZN(n3496) );
  and2 U3763 ( .A1(n3497), .A2(n3496), .Z(n3501) );
  inv1 U3764 ( .I(n3497), .ZN(n3499) );
  inv1 U3768 ( .I(n3503), .ZN(n3504) );
  or2 U3778 ( .A1(n3518), .A2(n2042), .Z(n3521) );
  or2 U3782 ( .A1(n3524), .A2(n2024), .Z(n3525) );
  and2 U3783 ( .A1(n3526), .A2(n3525), .Z(n3527) );
  or2 U3784 ( .A1(n3528), .A2(n3527), .Z(n3529) );
  and2 U3785 ( .A1(n3530), .A2(n3529), .Z(b11) );
  and2 U3786 ( .A1(n1919), .A2(n2028), .Z(n3534) );
  and2 U3787 ( .A1(n3532), .A2(n3531), .Z(n3533) );
  or2 U3788 ( .A1(n3534), .A2(n3533), .Z(n3536) );
  and2 U3789 ( .A1(n3535), .A2(n3536), .Z(n3540) );
  inv1 U3790 ( .I(n3536), .ZN(n3537) );
  and2 U3791 ( .A1(n3538), .A2(n3537), .Z(n3539) );
  or2 U3792 ( .A1(n3540), .A2(n3539), .Z(n3545) );
  inv1 U3793 ( .I(n3545), .ZN(n3547) );
  and2 U3794 ( .A1(n1454), .A2(n3547), .Z(n3543) );
  inv1 U3795 ( .I(n1454), .ZN(n3541) );
  and2 U3796 ( .A1(n3541), .A2(n3545), .Z(n3542) );
  or2 U3797 ( .A1(n3543), .A2(n3542), .Z(n3648) );
  inv1 U3798 ( .I(n3648), .ZN(n3544) );
  or2 U3799 ( .A1(n3544), .A2(n3647), .Z(n3574) );
  and2 U3800 ( .A1(n3546), .A2(n3545), .Z(n3550) );
  and2 U3801 ( .A1(n3548), .A2(n3547), .Z(n3549) );
  or2 U3802 ( .A1(n3550), .A2(n3549), .Z(n3567) );
  inv1 U3803 ( .I(n3555), .ZN(n3553) );
  inv1 U3804 ( .I(n3551), .ZN(n3552) );
  or2 U3805 ( .A1(n3553), .A2(n3552), .Z(n3557) );
  or2 U3806 ( .A1(n3555), .A2(n2949), .Z(n3556) );
  and2 U3807 ( .A1(n3557), .A2(n3556), .Z(n3558) );
  inv1 U3809 ( .I(n3562), .ZN(n3560) );
  inv1 U3813 ( .I(n3568), .ZN(n3566) );
  inv1 U3815 ( .I(n3567), .ZN(n3569) );
  inv1 U3818 ( .I(n3650), .ZN(n3572) );
  or2 U3823 ( .A1(n3577), .A2(n3576), .Z(n3582) );
  and2 U3824 ( .A1(n3579), .A2(n3578), .Z(n3580) );
  or2 U3825 ( .A1(n3580), .A2(n3625), .Z(n3583) );
  inv1 U3826 ( .I(n3583), .ZN(n3581) );
  and2 U3827 ( .A1(n3582), .A2(n3581), .Z(n3586) );
  inv1 U3828 ( .I(n3582), .ZN(n3584) );
  and2 U3829 ( .A1(n3584), .A2(n3583), .Z(n3585) );
  or2 U3830 ( .A1(n3586), .A2(n3585), .Z(n3588) );
  inv1 U3831 ( .I(n3588), .ZN(n3587) );
  and2 U3833 ( .A1(n3616), .A2(n3588), .Z(n3589) );
  and2 U3835 ( .A1(n3591), .A2(n3612), .Z(n3594) );
  and2 U3837 ( .A1(n3592), .A2(n3613), .Z(n3593) );
  and2 U3840 ( .A1(n3595), .A2(n2002), .Z(n3596) );
  or2 U3841 ( .A1(n3597), .A2(n3596), .Z(n3601) );
  inv1 U3842 ( .I(n3598), .ZN(n3599) );
  or2 U3843 ( .A1(n3599), .A2(n3617), .Z(n3602) );
  inv1 U3844 ( .I(n3602), .ZN(n3600) );
  and2 U3845 ( .A1(n3601), .A2(n3600), .Z(n3605) );
  inv1 U3846 ( .I(n3601), .ZN(n3603) );
  and2 U3847 ( .A1(n3603), .A2(n3602), .Z(n3604) );
  or2 U3848 ( .A1(n3605), .A2(n3604), .Z(n3608) );
  inv1 U3849 ( .I(n3608), .ZN(n3606) );
  or2 U3854 ( .A1(n3640), .A2(x6), .Z(n3637) );
  and2 U3855 ( .A1(n3625), .A2(n2057), .Z(n3615) );
  and2 U3857 ( .A1(n3616), .A2(n3620), .Z(n3618) );
  inv1 U3859 ( .I(n3621), .ZN(n3619) );
  and2 U3860 ( .A1(n3620), .A2(n3619), .Z(n3624) );
  inv1 U3861 ( .I(n3620), .ZN(n3622) );
  and2 U3862 ( .A1(n3622), .A2(n3621), .Z(n3623) );
  or2 U3864 ( .A1(n3626), .A2(n3625), .Z(n3629) );
  inv1 U3865 ( .I(n3629), .ZN(n3627) );
  or2 U3874 ( .A1(n3639), .A2(n3638), .Z(n3656) );
  inv1 U3877 ( .I(n3642), .ZN(n3644) );
  or2 U3880 ( .A1(n3648), .A2(n3647), .Z(n3652) );
  or2 U3881 ( .A1(n3650), .A2(n3649), .Z(n3651) );
  and2 U3882 ( .A1(n3652), .A2(n3651), .Z(n3653) );
  and2 U3884 ( .A1(n3656), .A2(n3655), .Z(c11) );
  inv1f U1956 ( .I(n2607), .ZN(n1989) );
  inv1f U1957 ( .I(n2091), .ZN(n2094) );
  inv1f U1959 ( .I(n2620), .ZN(n3062) );
  and2f U1963 ( .A1(n3420), .A2(n3148), .Z(n3151) );
  or2f U1964 ( .A1(n2142), .A2(n3420), .Z(n1986) );
  inv1 U1965 ( .I(n3420), .ZN(n3418) );
  or2f U1967 ( .A1(n2237), .A2(n1925), .Z(n2242) );
  inv1 U1968 ( .I(n3407), .ZN(n3409) );
  or2f U1971 ( .A1(n3023), .A2(n2995), .Z(n3407) );
  inv1f U1972 ( .I(n3401), .ZN(n3403) );
  or2f U1975 ( .A1(n3360), .A2(n3048), .Z(n1994) );
  inv1f U1977 ( .I(n2595), .ZN(n3048) );
  or2f U1979 ( .A1(n898), .A2(n3679), .Z(n897) );
  inv1 U1980 ( .I(n2983), .ZN(n2672) );
  or2f U1981 ( .A1(n1974), .A2(n1975), .Z(n2983) );
  or2 U1983 ( .A1(n3079), .A2(n3253), .Z(n2046) );
  or2f U1985 ( .A1(n3041), .A2(n3253), .Z(n3042) );
  or2f U1987 ( .A1(n2692), .A2(n3070), .Z(n3253) );
  and2f U1989 ( .A1(n3667), .A2(n2848), .Z(n2844) );
  or2f U1991 ( .A1(n2222), .A2(n2457), .Z(n2224) );
  and2f U1993 ( .A1(n2118), .A2(o), .Z(n1931) );
  inv1f U1994 ( .I(n2119), .ZN(n2106) );
  or2f U1995 ( .A1(n1915), .A2(n1919), .Z(n2960) );
  or2f U1998 ( .A1(n2134), .A2(n3134), .Z(n2137) );
  inv1f U1999 ( .I(n2132), .ZN(n3134) );
  inv1 U2000 ( .I(f), .ZN(n1930) );
  inv1f U2001 ( .I(n2419), .ZN(n2888) );
  or2f U2004 ( .A1(n2412), .A2(n2411), .Z(n2419) );
  and2f U2006 ( .A1(n2079), .A2(n3693), .Z(n1333) );
  inv1f U2007 ( .I(n2072), .ZN(n2079) );
  or2f U2010 ( .A1(n2649), .A2(n2648), .Z(n3218) );
  and2f U2014 ( .A1(n2068), .A2(n3217), .Z(n2649) );
  inv1f U2016 ( .I(n2029), .ZN(n3706) );
  inv1f U2022 ( .I(n3706), .ZN(n3707) );
  inv1f U2024 ( .I(n3706), .ZN(n3709) );
  inv1f U2027 ( .I(n3706), .ZN(n3708) );
  inv1f U2031 ( .I(n2261), .ZN(n2793) );
  or2f U2034 ( .A1(n2257), .A2(n2535), .Z(n2261) );
  inv1 U2037 ( .I(f), .ZN(n3710) );
  inv1 U2038 ( .I(f), .ZN(n2120) );
  inv1 U2039 ( .I(f), .ZN(n2122) );
  inv1f U2040 ( .I(f), .ZN(n1951) );
  inv1f U2042 ( .I(f), .ZN(n2118) );
  inv1f U2046 ( .I(f), .ZN(n1946) );
  inv1 U2047 ( .I(n2079), .ZN(n1944) );
  inv1f U2048 ( .I(f), .ZN(n1928) );
  or2f U2049 ( .A1(n2472), .A2(n3707), .Z(n2594) );
  or2f U2050 ( .A1(n2478), .A2(n3708), .Z(n2590) );
  or2f U2051 ( .A1(n2480), .A2(n3709), .Z(n2591) );
  or2f U2052 ( .A1(n2480), .A2(n3707), .Z(n1992) );
  inv1f U2054 ( .I(n3708), .ZN(n2101) );
  and2 U2057 ( .A1(i1), .A2(n2817), .Z(n2240) );
  and2 U2063 ( .A1(n2444), .A2(n2080), .Z(n2445) );
  or2 U2064 ( .A1(n2841), .A2(n2842), .Z(n2840) );
  and2 U2065 ( .A1(r3), .A2(f), .Z(n2257) );
  and2 U2066 ( .A1(n3358), .A2(n3314), .Z(n3315) );
  or2 U2067 ( .A1(n2341), .A2(n2340), .Z(n2352) );
  or2 U2069 ( .A1(n2248), .A2(n2247), .Z(n960) );
  and2 U2070 ( .A1(f), .A2(n2246), .Z(n2247) );
  and2 U2071 ( .A1(g3), .A2(f), .Z(n2237) );
  or2 U2072 ( .A1(n2770), .A2(n2771), .Z(n2769) );
  inv1 U2078 ( .I(n3172), .ZN(n3174) );
  and2 U2081 ( .A1(n900), .A2(n901), .Z(n898) );
  and2 U2084 ( .A1(n1011), .A2(n1012), .Z(n1009) );
  and2 U2086 ( .A1(n1928), .A2(j), .Z(n1962) );
  and2 U2089 ( .A1(n3358), .A2(n3370), .Z(n2706) );
  inv1 U2091 ( .I(n3178), .ZN(n3179) );
  inv1 U2092 ( .I(n3373), .ZN(n3375) );
  or2 U2093 ( .A1(n3326), .A2(n3325), .Z(n3327) );
  or2 U2094 ( .A1(n684), .A2(n685), .Z(n682) );
  or2 U2098 ( .A1(n630), .A2(n631), .Z(n628) );
  or2 U2099 ( .A1(n3314), .A2(n3308), .Z(n3026) );
  or2 U2104 ( .A1(n2447), .A2(n3707), .Z(n2687) );
  or2 U2105 ( .A1(n2653), .A2(n2652), .Z(n3079) );
  and2 U2111 ( .A1(n3462), .A2(n3486), .Z(n3465) );
  and2 U2113 ( .A1(n3502), .A2(n3503), .Z(n3507) );
  and2 U2114 ( .A1(n3486), .A2(n3485), .Z(n3489) );
  inv1 U2120 ( .I(n2970), .ZN(n2969) );
  or2 U2121 ( .A1(n2573), .A2(n2572), .Z(n2574) );
  and2 U2123 ( .A1(n2571), .A2(n2570), .Z(n2572) );
  inv1 U2124 ( .I(n2468), .ZN(n3663) );
  inv1 U2125 ( .I(n2373), .ZN(n3673) );
  or2 U2126 ( .A1(n2295), .A2(n2294), .Z(n888) );
  and2 U2130 ( .A1(n2292), .A2(n2293), .Z(n2295) );
  or2 U2131 ( .A1(n2226), .A2(n2225), .Z(n999) );
  or2 U2132 ( .A1(n3348), .A2(n3323), .Z(n3314) );
  and2 U2134 ( .A1(n2432), .A2(f), .Z(n2433) );
  or2 U2135 ( .A1(n2647), .A2(n2646), .Z(n3217) );
  inv1 U2136 ( .I(n3026), .ZN(n3371) );
  or2 U2137 ( .A1(n2680), .A2(n2679), .Z(n3255) );
  or2 U2140 ( .A1(n3555), .A2(n3554), .Z(n2618) );
  inv1 U2143 ( .I(n3113), .ZN(n3120) );
  inv1 U2147 ( .I(n3273), .ZN(n3292) );
  or2 U2148 ( .A1(n3266), .A2(n3268), .Z(n3267) );
  and2 U2150 ( .A1(n3569), .A2(n3568), .Z(n3570) );
  and2 U2153 ( .A1(n3607), .A2(n3606), .Z(n3611) );
  and2 U2155 ( .A1(n2885), .A2(n2884), .Z(n2906) );
  or2 U2156 ( .A1(n2987), .A2(n2986), .Z(n2988) );
  or2 U2157 ( .A1(n2828), .A2(n2827), .Z(n2829) );
  inv1 U2158 ( .I(n3189), .ZN(n3190) );
  or2 U2159 ( .A1(n2594), .A2(b1), .Z(n2595) );
  or2 U2160 ( .A1(n1918), .A2(n2053), .Z(n2051) );
  inv1 U2161 ( .I(n2024), .ZN(n3522) );
  or2 U2162 ( .A1(n1990), .A2(n3409), .Z(n3411) );
  or2 U2164 ( .A1(n3408), .A2(n3407), .Z(n3412) );
  inv1 U2166 ( .I(n3518), .ZN(n3481) );
  or2 U2168 ( .A1(n512), .A2(n513), .Z(n395) );
  or2 U2175 ( .A1(n618), .A2(n619), .Z(n617) );
  or2 U2176 ( .A1(n846), .A2(n847), .Z(s9) );
  inv1 U2178 ( .I(n3301), .ZN(n3302) );
  inv1 U2180 ( .I(n2094), .ZN(n2002) );
  inv1f U2181 ( .I(n2127), .ZN(n2141) );
  inv1f U2184 ( .I(n767), .ZN(n3677) );
  inv1f U2188 ( .I(n2917), .ZN(n3625) );
  and2f U2189 ( .A1(n3710), .A2(l1), .Z(n1950) );
  and2f U2190 ( .A1(n2111), .A2(i), .Z(n1949) );
  inv1f U2191 ( .I(n2059), .ZN(n2061) );
  or2f U2192 ( .A1(n2845), .A2(n2895), .Z(n2847) );
  inv1f U2193 ( .I(n3463), .ZN(n3462) );
  or2 U2194 ( .A1(n3183), .A2(n3186), .Z(n3169) );
  or2f U2195 ( .A1(n2639), .A2(n2646), .Z(n3186) );
  or2f U2196 ( .A1(n3065), .A2(n2010), .Z(n3081) );
  or2f U2197 ( .A1(n2151), .A2(n1924), .Z(n1920) );
  or2f U2198 ( .A1(n2161), .A2(n2619), .Z(n3554) );
  and2f U2199 ( .A1(n2069), .A2(n2641), .Z(n2068) );
  and2 U2200 ( .A1(n1981), .A2(n2056), .Z(n3577) );
  or2f U2201 ( .A1(n2656), .A2(n2017), .Z(n2056) );
  and2f U2202 ( .A1(c), .A2(d), .Z(n2029) );
  inv1 U2204 ( .I(n2101), .ZN(n2104) );
  or2f U2205 ( .A1(n2660), .A2(h6), .Z(n2664) );
  or2f U2206 ( .A1(n2623), .A2(n3139), .Z(n2979) );
  or2f U2207 ( .A1(n2136), .A2(n2696), .Z(n3139) );
  or2f U2208 ( .A1(n2674), .A2(n3132), .Z(n3446) );
  and2f U2209 ( .A1(n1982), .A2(n2655), .Z(n1981) );
  and2f U2218 ( .A1(n2507), .A2(n2169), .Z(n1983) );
  and2 U2223 ( .A1(e5), .A2(f), .Z(n2569) );
  and2 U2224 ( .A1(c5), .A2(f), .Z(n2563) );
  and2 U2225 ( .A1(n1988), .A2(n3441), .Z(n3444) );
  and2f U2226 ( .A1(n1989), .A2(n2606), .Z(n1988) );
  or2f U2236 ( .A1(n2066), .A2(n3446), .Z(n3115) );
  and2f U2237 ( .A1(n3446), .A2(n3445), .Z(n3450) );
  inv1f U2238 ( .I(n3446), .ZN(n3448) );
  or2f U2239 ( .A1(n2559), .A2(l6), .Z(n2157) );
  inv1f U2240 ( .I(n2557), .ZN(n2559) );
  or2 U2247 ( .A1(n2945), .A2(n1919), .Z(n3555) );
  and2f U2252 ( .A1(n2842), .A2(n2841), .Z(n2843) );
  inv1f U2270 ( .I(n2224), .ZN(n2842) );
  inv1f U2271 ( .I(n2157), .ZN(n2947) );
  inv1f U2280 ( .I(f), .ZN(n2119) );
  inv1f U2282 ( .I(f), .ZN(n2049) );
  or2 U2283 ( .A1(n2323), .A2(n2322), .Z(n767) );
  or2 U2288 ( .A1(n2888), .A2(t5), .Z(n2417) );
  and2 U2289 ( .A1(b4), .A2(n2793), .Z(n2259) );
  and2 U2291 ( .A1(n2840), .A2(n2839), .Z(n2845) );
  and2 U2292 ( .A1(n3184), .A2(n3183), .Z(n3188) );
  and2 U2293 ( .A1(n3191), .A2(n3190), .Z(n3192) );
  and2 U2300 ( .A1(n2687), .A2(n2450), .Z(n2452) );
  or2 U2405 ( .A1(n2216), .A2(n2215), .Z(n2217) );
  and2 U2406 ( .A1(n2633), .A2(n2108), .Z(n2412) );
  or2 U2415 ( .A1(n3493), .A2(n3442), .Z(n3482) );
  or2 U2418 ( .A1(n2156), .A2(n1950), .Z(n2557) );
  and2 U2423 ( .A1(n635), .A2(n636), .Z(n633) );
  inv1 U2425 ( .I(n637), .ZN(n636) );
  and2 U2426 ( .A1(n2866), .A2(n2865), .Z(n2869) );
  or2 U2427 ( .A1(n2864), .A2(n2894), .Z(n2865) );
  and2 U2444 ( .A1(n2859), .A2(n2858), .Z(n2864) );
  or2 U2445 ( .A1(n2844), .A2(n2843), .Z(n2895) );
  and2 U2447 ( .A1(n2771), .A2(n2770), .Z(n2772) );
  or2 U2456 ( .A1(n2816), .A2(n2817), .Z(n2731) );
  inv1 U2457 ( .I(n3064), .ZN(n2048) );
  and2 U2467 ( .A1(n3172), .A2(n3171), .Z(n3176) );
  or2 U2468 ( .A1(n3166), .A2(n3218), .Z(n1963) );
  or2 U2470 ( .A1(n3204), .A2(n3203), .Z(n3228) );
  inv1 U2474 ( .I(n3228), .ZN(n3229) );
  or2 U2476 ( .A1(n3461), .A2(n3460), .Z(n3486) );
  inv1 U2477 ( .I(n3486), .ZN(n3487) );
  inv1 U2509 ( .I(n1969), .ZN(n2570) );
  or2 U2525 ( .A1(n740), .A2(n741), .Z(n737) );
  or2 U2528 ( .A1(n744), .A2(n742), .Z(n745) );
  and2 U2567 ( .A1(n1010), .A2(n1009), .Z(n1006) );
  or2 U2569 ( .A1(n895), .A2(n896), .Z(n893) );
  inv1 U2570 ( .I(n3180), .ZN(n3177) );
  or2 U2595 ( .A1(n2697), .A2(n2696), .Z(n2986) );
  and2 U2635 ( .A1(n2985), .A2(n2984), .Z(n2987) );
  or2 U2636 ( .A1(n2078), .A2(n3132), .Z(n2984) );
  or2 U2637 ( .A1(n2671), .A2(n3575), .Z(n2942) );
  inv1 U2701 ( .I(n3350), .ZN(n3348) );
  inv1 U2703 ( .I(n2687), .ZN(n2675) );
  or2 U2704 ( .A1(n2431), .A2(n3709), .Z(n2579) );
  and2 U2710 ( .A1(s4), .A2(f), .Z(n2529) );
  or2 U2724 ( .A1(n2044), .A2(u6), .Z(n2127) );
  or2 U2727 ( .A1(n2124), .A2(n1947), .Z(n2507) );
  or2 U2730 ( .A1(n3613), .A2(n3614), .Z(n1954) );
  inv1 U2731 ( .I(n3607), .ZN(n3609) );
  inv1 U2749 ( .I(n3614), .ZN(n1968) );
  inv1 U2750 ( .I(n2664), .ZN(n3617) );
  and2 U2753 ( .A1(n2570), .A2(n2018), .Z(n2017) );
  inv1 U2758 ( .I(n681), .ZN(n680) );
  or2 U2759 ( .A1(n2429), .A2(n2428), .Z(n623) );
  inv1 U2782 ( .I(n2254), .ZN(n3703) );
  or2 U2788 ( .A1(n2879), .A2(n2878), .Z(n2880) );
  inv1 U2797 ( .I(n2877), .ZN(n2878) );
  and2 U2800 ( .A1(n2901), .A2(n2900), .Z(n2902) );
  and2 U2849 ( .A1(n2887), .A2(n2886), .Z(n2901) );
  inv1 U2858 ( .I(n2999), .ZN(n3008) );
  and2 U2864 ( .A1(n2015), .A2(n2633), .Z(n2014) );
  or2 U2893 ( .A1(n2705), .A2(n2704), .Z(n3370) );
  inv1 U2900 ( .I(n3253), .ZN(n3256) );
  or2 U2903 ( .A1(n3502), .A2(n3462), .Z(n3447) );
  and2 U2904 ( .A1(n2061), .A2(n3234), .Z(n3239) );
  or2 U2919 ( .A1(n3233), .A2(n3235), .Z(n3234) );
  or2 U2922 ( .A1(n3290), .A2(n3293), .Z(n3291) );
  inv1 U2923 ( .I(n3510), .ZN(n3508) );
  and2 U2937 ( .A1(n3509), .A2(n2042), .Z(n2006) );
  inv1 U2940 ( .I(n2042), .ZN(n2060) );
  inv1 U2945 ( .I(n3509), .ZN(n3511) );
  and2 U2947 ( .A1(n3478), .A2(n3477), .Z(n3479) );
  inv1 U2948 ( .I(n1981), .ZN(n3575) );
  inv1 U2964 ( .I(n2070), .ZN(n3578) );
  or2 U2968 ( .A1(n557), .A2(n3663), .Z(n553) );
  or2 U2969 ( .A1(n888), .A2(n889), .Z(n887) );
  inv1 U2970 ( .I(n3183), .ZN(n3185) );
  or2 U2975 ( .A1(n2035), .A2(n2036), .Z(n2034) );
  inv1 U2976 ( .I(n1988), .ZN(n3442) );
  inv1 U2977 ( .I(n2611), .ZN(n2022) );
  or2 U2980 ( .A1(n3384), .A2(n3409), .Z(n3385) );
  or2 U2983 ( .A1(n3346), .A2(n3407), .Z(n3386) );
  or2 U2985 ( .A1(n3572), .A2(n3649), .Z(n3573) );
  or2 U2987 ( .A1(n3641), .A2(x6), .Z(n3646) );
  inv1 U2989 ( .I(n3640), .ZN(n3641) );
  or2 U2990 ( .A1(n728), .A2(n729), .Z(n616) );
  or2 U2991 ( .A1(n730), .A2(n731), .Z(n729) );
  or2 U2995 ( .A1(n1956), .A2(n1957), .Z(t9) );
  and2 U3001 ( .A1(n3189), .A2(n3001), .Z(n3004) );
  inv1 U3002 ( .I(n2082), .ZN(n3049) );
  and2 U3007 ( .A1(n3659), .A2(n3083), .Z(n3086) );
  or2 U3008 ( .A1(n3083), .A2(n3659), .Z(n3084) );
  and2 U3015 ( .A1(n3089), .A2(n3088), .Z(n3094) );
  inv1 U3016 ( .I(n3303), .ZN(n3300) );
  and2 U3017 ( .A1(n3515), .A2(n3514), .Z(n3516) );
  or2 U3018 ( .A1(n3079), .A2(n3253), .Z(n2698) );
  inv1 U3022 ( .I(n3341), .ZN(n3343) );
  and2f U3026 ( .A1(n3341), .A2(n3340), .Z(n3345) );
  and2f U3027 ( .A1(n3320), .A2(n3319), .Z(n3321) );
  inv1 U3033 ( .I(n902), .ZN(n901) );
  and2 U3035 ( .A1(n3679), .A2(n898), .Z(n895) );
  and2f U3036 ( .A1(n903), .A2(n904), .Z(n902) );
  or2f U3039 ( .A1(n2823), .A2(n1961), .Z(n1959) );
  or2 U3040 ( .A1(n1918), .A2(n3313), .Z(n1917) );
  or2f U3041 ( .A1(n3400), .A2(n3401), .Z(n3397) );
  inv1 U3042 ( .I(n2096), .ZN(n3396) );
  and2f U3043 ( .A1(n2072), .A2(p), .Z(n1952) );
  or2f U3045 ( .A1(n3513), .A2(n3512), .Z(n3519) );
  inv1 U3049 ( .I(n1004), .ZN(n2223) );
  and2f U3050 ( .A1(n996), .A2(n997), .Z(n940) );
  or2f U3057 ( .A1(n2533), .A2(n2532), .Z(n2534) );
  or2f U3059 ( .A1(n3654), .A2(n3653), .Z(n3655) );
  and2 U3060 ( .A1(n3626), .A2(n2094), .Z(n3597) );
  and2f U3064 ( .A1(n1910), .A2(n2039), .Z(n2989) );
  or2f U3065 ( .A1(n1911), .A2(n2983), .Z(n1910) );
  inv1 U3068 ( .I(n1910), .ZN(n2041) );
  inv1 U3069 ( .I(n555), .ZN(n554) );
  and2f U3074 ( .A1(n3663), .A2(n557), .Z(n555) );
  or2f U3075 ( .A1(n2433), .A2(n3709), .Z(n2627) );
  and2f U3076 ( .A1(n2023), .A2(n3371), .Z(n3045) );
  or2f U3082 ( .A1(n3456), .A2(n3455), .Z(n3459) );
  or2f U3083 ( .A1(n3465), .A2(n3464), .Z(n3476) );
  or2f U3087 ( .A1(n3523), .A2(n3522), .Z(n3526) );
  or2f U3092 ( .A1(n3383), .A2(n3382), .Z(n1990) );
  and2f U3093 ( .A1(n2904), .A2(n2903), .Z(n2905) );
  and2f U3094 ( .A1(n2856), .A2(n2855), .Z(n2859) );
  and2f U3100 ( .A1(n3404), .A2(n3401), .Z(n2096) );
  or2f U3101 ( .A1(n2445), .A2(n3708), .Z(n2678) );
  or2f U3123 ( .A1(n3060), .A2(n2981), .Z(n1971) );
  or2f U3157 ( .A1(n2004), .A2(n2005), .Z(n2003) );
  and2f U3161 ( .A1(n1988), .A2(n3494), .Z(n2615) );
  and2f U3191 ( .A1(n1988), .A2(n1995), .Z(n2077) );
  and2 U3193 ( .A1(t4), .A2(f), .Z(n2523) );
  or2f U3201 ( .A1(n616), .A2(n617), .Z(r9) );
  or2f U3203 ( .A1(n746), .A2(n747), .Z(n742) );
  or2f U3204 ( .A1(n3594), .A2(n3593), .Z(n3607) );
  or2f U3205 ( .A1(n3082), .A2(n3274), .Z(n3083) );
  and2f U3206 ( .A1(n3081), .A2(n3080), .Z(n3082) );
  or2f U3207 ( .A1(n3199), .A2(n3198), .Z(n3202) );
  or2f U3217 ( .A1(n3232), .A2(n3231), .Z(n3235) );
  and2f U3219 ( .A1(n3230), .A2(n3229), .Z(n3231) );
  and2f U3223 ( .A1(n3630), .A2(n3629), .Z(n3631) );
  inv1f U3224 ( .I(n3628), .ZN(n3630) );
  or2f U3227 ( .A1(n2060), .A2(n3493), .Z(n3113) );
  and2f U3232 ( .A1(n2065), .A2(n2655), .Z(n1987) );
  or2f U3234 ( .A1(n3399), .A2(n3398), .Z(n3416) );
  and2f U3235 ( .A1(n410), .A2(n411), .Z(n406) );
  or2f U3236 ( .A1(n2830), .A2(n2998), .Z(n2879) );
  inv1f U3239 ( .I(n1998), .ZN(n3635) );
  or2f U3241 ( .A1(n1999), .A2(n2000), .Z(n1998) );
  and2f U3248 ( .A1(n2626), .A2(n2625), .Z(n2644) );
  and2f U3250 ( .A1(n2143), .A2(n3418), .Z(n2134) );
  or2f U3256 ( .A1(n3020), .A2(n3022), .Z(n2995) );
  or2f U3323 ( .A1(n3036), .A2(n3035), .Z(c10) );
  or2f U3324 ( .A1(n3023), .A2(n3022), .Z(n3024) );
  or2f U3325 ( .A1(n3062), .A2(n3060), .Z(n2982) );
  or2f U3327 ( .A1(n3554), .A2(n2157), .Z(n2085) );
  or2f U3330 ( .A1(n3023), .A2(n3020), .Z(n3044) );
  or2f U3331 ( .A1(n2619), .A2(n1919), .Z(n2073) );
  or2f U3332 ( .A1(n3501), .A2(n3500), .Z(n3503) );
  and2f U3333 ( .A1(n3499), .A2(n3498), .Z(n3500) );
  or2f U3334 ( .A1(n2613), .A2(n2612), .Z(n3494) );
  and2f U3335 ( .A1(n3574), .A2(n3573), .Z(n3639) );
  and2f U3341 ( .A1(n3563), .A2(n3562), .Z(n3564) );
  or2f U3342 ( .A1(n3559), .A2(n3558), .Z(n3562) );
  inv1f U3343 ( .I(n2547), .ZN(n2549) );
  or2f U3344 ( .A1(n1945), .A2(n2152), .Z(n2547) );
  or2f U3346 ( .A1(n3383), .A2(n3382), .Z(n3410) );
  or2f U3367 ( .A1(n3363), .A2(n3362), .Z(n3366) );
  and2f U3369 ( .A1(n3361), .A2(n3365), .Z(n3363) );
  or2f U3373 ( .A1(n848), .A2(n849), .Z(n847) );
  and2f U3374 ( .A1(n3189), .A2(n3167), .Z(n2092) );
  and2f U3379 ( .A1(n3040), .A2(n3039), .Z(n3041) );
  and2f U3381 ( .A1(n3038), .A2(n2047), .Z(n3040) );
  and2f U3383 ( .A1(n1917), .A2(n2083), .Z(n2082) );
  or2f U3384 ( .A1(n2671), .A2(n3575), .Z(n2065) );
  and2f U3387 ( .A1(n3575), .A2(n2057), .Z(n3576) );
  or2f U3388 ( .A1(n940), .A2(n941), .Z(n846) );
  and2 U3389 ( .A1(n946), .A2(n945), .Z(n942) );
  or2f U3402 ( .A1(n2582), .A2(f), .Z(n3614) );
  and2f U3420 ( .A1(n2068), .A2(n3008), .Z(n3000) );
  or2f U3422 ( .A1(n2616), .A2(n3491), .Z(n2078) );
  or2f U3423 ( .A1(n2075), .A2(n2076), .Z(n2616) );
  and2f U3424 ( .A1(n3561), .A2(n3560), .Z(n3565) );
  and2f U3427 ( .A1(n1923), .A2(n3587), .Z(n3590) );
  or2f U3429 ( .A1(n3618), .A2(n3617), .Z(n3621) );
  or2f U3438 ( .A1(n2917), .A2(n1923), .Z(n2662) );
  and2f U3443 ( .A1(n2059), .A2(n3210), .Z(n3215) );
  or2f U3459 ( .A1(n3209), .A2(n3212), .Z(n3210) );
  or2f U3460 ( .A1(n3176), .A2(n3175), .Z(n3178) );
  and2f U3463 ( .A1(n2067), .A2(n2645), .Z(n2647) );
  and2f U3465 ( .A1(n2912), .A2(n2880), .Z(n2885) );
  or2f U3492 ( .A1(n2875), .A2(n2890), .Z(n2887) );
  or2f U3508 ( .A1(n3023), .A2(n3020), .Z(n2023) );
  or2f U3514 ( .A1(n3538), .A2(n3531), .Z(n2945) );
  and2f U3515 ( .A1(n3292), .A2(n3291), .Z(n3297) );
  and2f U3517 ( .A1(n3287), .A2(n3286), .Z(n3288) );
  and2f U3519 ( .A1(a6), .A2(n2689), .Z(n2680) );
  inv1f U3520 ( .I(n2003), .ZN(n3514) );
  and2f U3523 ( .A1(n2042), .A2(n3512), .Z(n2005) );
  or2f U3527 ( .A1(r9), .A2(r8), .Z(n612) );
  or2f U3533 ( .A1(n3674), .A2(n3673), .Z(n734) );
  and2f U3537 ( .A1(n1980), .A2(n3633), .Z(n3634) );
  or2f U3540 ( .A1(n1980), .A2(n3632), .Z(n2000) );
  and2f U3543 ( .A1(n3406), .A2(n3405), .Z(n3414) );
  or2f U3544 ( .A1(n3404), .A2(n3403), .Z(n3405) );
  or2f U3545 ( .A1(n1915), .A2(n2086), .Z(n2084) );
  and2f U3558 ( .A1(n2701), .A2(n2700), .Z(n2711) );
  and2f U3559 ( .A1(n3273), .A2(n3267), .Z(n3272) );
  and2f U3560 ( .A1(n3120), .A2(n2037), .Z(n2035) );
  or2f U3561 ( .A1(n3177), .A2(n2014), .Z(n3183) );
  and2f U3565 ( .A1(n3509), .A2(n3508), .Z(n3513) );
  and2f U3566 ( .A1(n3521), .A2(n3520), .Z(n3528) );
  or2f U3588 ( .A1(n3519), .A2(n2060), .Z(n3520) );
  or2f U3589 ( .A1(n3409), .A2(n3314), .Z(n3053) );
  inv1f U3592 ( .I(n3255), .ZN(n3252) );
  inv1f U3593 ( .I(n3380), .ZN(n3378) );
  and2f U3601 ( .A1(n3373), .A2(n3372), .Z(n3377) );
  or2f U3602 ( .A1(n3369), .A2(n3368), .Z(n3373) );
  or2f U3603 ( .A1(n677), .A2(n678), .Z(n676) );
  and2f U3604 ( .A1(n679), .A2(n680), .Z(n677) );
  and2f U3607 ( .A1(n682), .A2(n683), .Z(n681) );
  and2f U3608 ( .A1(n2906), .A2(n1958), .Z(n1956) );
  inv1f U3610 ( .I(n2213), .ZN(n2889) );
  or2f U3612 ( .A1(n2208), .A2(n1921), .Z(n2213) );
  or2f U3617 ( .A1(n1009), .A2(n1010), .Z(n1008) );
  or2f U3620 ( .A1(n1006), .A2(n1007), .Z(n1004) );
  and2 U3622 ( .A1(n1004), .A2(n2842), .Z(n2225) );
  or2f U3623 ( .A1(n3635), .A2(n3634), .Z(n2001) );
  or2f U3626 ( .A1(n3635), .A2(n3634), .Z(n3642) );
  or2f U3627 ( .A1(n3632), .A2(n3631), .Z(n3633) );
  and2f U3642 ( .A1(n2057), .A2(n3626), .Z(n2667) );
  and2f U3643 ( .A1(n3324), .A2(n3349), .Z(n3325) );
  or2f U3644 ( .A1(n3345), .A2(n3344), .Z(n3408) );
  and2f U3645 ( .A1(n3343), .A2(n3342), .Z(n3344) );
  or2f U3647 ( .A1(n3322), .A2(n3321), .Z(n3347) );
  and2f U3653 ( .A1(n3318), .A2(n3317), .Z(n3322) );
  or2f U3654 ( .A1(n3480), .A2(n3479), .Z(n3518) );
  inv1f U3655 ( .I(n2118), .ZN(n2080) );
  inv1f U3656 ( .I(n2978), .ZN(n3132) );
  or2f U3657 ( .A1(n623), .A2(n624), .Z(n622) );
  inv1f U3662 ( .I(n632), .ZN(n631) );
  and2f U3665 ( .A1(n3462), .A2(n2021), .Z(n2613) );
  and2f U3666 ( .A1(n950), .A2(n2733), .Z(n2254) );
  or2f U3667 ( .A1(n945), .A2(n946), .Z(n944) );
  and2f U3668 ( .A1(n947), .A2(n3703), .Z(n945) );
  or2f U3669 ( .A1(n3565), .A2(n3564), .Z(n3568) );
  or2f U3670 ( .A1(n3571), .A2(n3570), .Z(n3650) );
  and2f U3672 ( .A1(n3567), .A2(n3566), .Z(n3571) );
  and2f U3673 ( .A1(n1951), .A2(m1), .Z(n1945) );
  and2f U3675 ( .A1(n1916), .A2(n2153), .Z(n1915) );
  inv1f U3676 ( .I(n2155), .ZN(n1916) );
  or2f U3681 ( .A1(n2869), .A2(n2891), .Z(n2872) );
  and2f U3686 ( .A1(n3412), .A2(n3411), .Z(n3413) );
  and2f U3689 ( .A1(n3375), .A2(n3374), .Z(n3376) );
  and2f U3690 ( .A1(n3323), .A2(n3306), .Z(n2704) );
  or2f U3691 ( .A1(n3578), .A2(n3579), .Z(n2917) );
  or2f U3692 ( .A1(n1968), .A2(n3591), .Z(n3579) );
  inv1f U3693 ( .I(n3592), .ZN(n3591) );
  and2f U3717 ( .A1(n3131), .A2(n2978), .Z(n2024) );
  and2f U3720 ( .A1(n1976), .A2(n1977), .Z(n3131) );
  or2f U3727 ( .A1(n3516), .A2(n3517), .Z(n3530) );
  and2f U3731 ( .A1(n3487), .A2(n2007), .Z(n3488) );
  and2f U3732 ( .A1(n3463), .A2(n3487), .Z(n3464) );
  and2f U3733 ( .A1(n3180), .A2(n3179), .Z(n3181) );
  or2f U3734 ( .A1(n3241), .A2(n3240), .Z(n3303) );
  and2f U3735 ( .A1(n3215), .A2(n3214), .Z(n3241) );
  or2f U3748 ( .A1(n3362), .A2(n3032), .Z(n3034) );
  and2f U3749 ( .A1(n3031), .A2(n3030), .Z(n3032) );
  and2f U3750 ( .A1(n2994), .A2(n2694), .Z(n3022) );
  and2f U3755 ( .A1(n2991), .A2(n2992), .Z(n2994) );
  or2f U3756 ( .A1(n2128), .A2(n2141), .Z(n2143) );
  and2f U3765 ( .A1(n1983), .A2(n2140), .Z(n2128) );
  or2f U3766 ( .A1(n2095), .A2(n3167), .Z(n3002) );
  and2f U3767 ( .A1(n3005), .A2(n2019), .Z(n2095) );
  or2f U3769 ( .A1(n2989), .A2(n2988), .Z(n2059) );
  or2f U3770 ( .A1(n2145), .A2(n3417), .Z(n2623) );
  or2f U3771 ( .A1(n1986), .A2(n2141), .Z(n2145) );
  or2f U3772 ( .A1(n2133), .A2(n3134), .Z(n3420) );
  inv1f U3773 ( .I(n3612), .ZN(n3613) );
  or2f U3774 ( .A1(n3590), .A2(n3589), .Z(n3612) );
  or2f U3775 ( .A1(n3611), .A2(n3610), .Z(n3640) );
  and2f U3776 ( .A1(n3609), .A2(n3608), .Z(n3610) );
  inv1f U3777 ( .I(f), .ZN(n2111) );
  or2f U3779 ( .A1(n2372), .A2(n2371), .Z(n2373) );
  and2f U3780 ( .A1(n2370), .A2(n2369), .Z(n2371) );
  and2f U3781 ( .A1(n2321), .A2(f), .Z(n2323) );
  or2f U3808 ( .A1(n2711), .A2(n2710), .Z(n2712) );
  and2f U3810 ( .A1(n2011), .A2(n2012), .Z(n2653) );
  and2f U3811 ( .A1(n2020), .A2(n2631), .Z(n2019) );
  and2f U3812 ( .A1(n999), .A2(n1000), .Z(n998) );
  inv1f U3814 ( .I(n2049), .ZN(n2108) );
  inv1f U3816 ( .I(n897), .ZN(n896) );
  or2f U3817 ( .A1(n3357), .A2(n3356), .Z(n3379) );
  and2f U3819 ( .A1(n3355), .A2(n3354), .Z(n3356) );
  and2f U3820 ( .A1(n3381), .A2(n3380), .Z(n3382) );
  or2f U3821 ( .A1(n3377), .A2(n3376), .Z(n3380) );
  and2f U3822 ( .A1(n3087), .A2(n2062), .Z(n3089) );
  and2f U3832 ( .A1(n3598), .A2(n2668), .Z(n2671) );
  or2f U3834 ( .A1(n2094), .A2(n1923), .Z(n3598) );
  and2f U3836 ( .A1(n3081), .A2(n3243), .Z(n2062) );
  or2f U3838 ( .A1(n2661), .A2(n3617), .Z(n1923) );
  or2f U3839 ( .A1(n3047), .A2(n3046), .Z(n3051) );
  or2f U3850 ( .A1(n3045), .A2(n3370), .Z(n3046) );
  inv1f U3851 ( .I(n2686), .ZN(n3023) );
  or2f U3852 ( .A1(n2685), .A2(n2684), .Z(n2686) );
  or2f U3853 ( .A1(n2158), .A2(n2947), .Z(n1919) );
  and2f U3856 ( .A1(n3637), .A2(n3636), .Z(n3638) );
  or2f U3858 ( .A1(n2001), .A2(n3643), .Z(n3636) );
  and2f U3863 ( .A1(n3628), .A2(n3627), .Z(n3632) );
  or2f U3866 ( .A1(n3624), .A2(n3623), .Z(n3628) );
  or2f U3867 ( .A1(n3615), .A2(n2002), .Z(n3620) );
  or2f U3868 ( .A1(n3299), .A2(n3298), .Z(n3301) );
  and2f U3869 ( .A1(n3272), .A2(n3271), .Z(n3299) );
  and2f U3870 ( .A1(n3297), .A2(n3296), .Z(n3298) );
  or2f U3871 ( .A1(n3289), .A2(n3288), .Z(n3293) );
  and2f U3872 ( .A1(n3659), .A2(n3248), .Z(n2692) );
  and2f U3873 ( .A1(n3305), .A2(n3304), .Z(z10) );
  or2f U3875 ( .A1(n3000), .A2(n3218), .Z(n3005) );
  or2f U3876 ( .A1(n3166), .A2(n3218), .Z(n3206) );
  or2f U3878 ( .A1(n3507), .A2(n3506), .Z(n3510) );
  and2f U3879 ( .A1(n3505), .A2(n3504), .Z(n3506) );
  and2f U3883 ( .A1(n3511), .A2(n3510), .Z(n3512) );
  and2f U3885 ( .A1(n2022), .A2(n2610), .Z(n2021) );
  inv1f U3886 ( .I(f), .ZN(n2072) );
  and2f U3887 ( .A1(n3386), .A2(n3385), .Z(n3399) );
  and2f U3888 ( .A1(n3379), .A2(n3378), .Z(n3383) );
  and2f U3889 ( .A1(n3358), .A2(n3371), .Z(n3360) );
  and2f U3890 ( .A1(n3646), .A2(n3645), .Z(n3654) );
  or2f U3891 ( .A1(n3644), .A2(n3643), .Z(n3645) );
  and2f U3892 ( .A1(n1954), .A2(n1967), .Z(n1980) );
  inv1f U3893 ( .I(n1928), .ZN(n2107) );
  or2f U3894 ( .A1(n2048), .A2(n3079), .Z(n2047) );
  and2f U3895 ( .A1(n2979), .A2(n2624), .Z(n2626) );
  or2f U3896 ( .A1(n2138), .A2(n3139), .Z(n2624) );
  or2f U3897 ( .A1(n2713), .A2(n2712), .Z(n3401) );
  and2f U3898 ( .A1(n3044), .A2(n2063), .Z(n2713) );
  or2f U3899 ( .A1(n3099), .A2(n2026), .Z(n2042) );
  or2f U3900 ( .A1(n2666), .A2(n2665), .Z(n3626) );
  and2f U3901 ( .A1(n3591), .A2(n2087), .Z(n2666) );
  and2f U3902 ( .A1(n3098), .A2(n3647), .Z(n3099) );
  inv1f U3903 ( .I(n1987), .ZN(n3647) );
endmodule

