
module C3540_iscas ( x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, 
        j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, 
        p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, t1, s1, r1, q1, p1, o1, 
        n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0 );
  input x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0,
         f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l,
         k, j, i, h, g, f, e, d, c, b, a;
  output t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1,
         c1, b1, a1, z0, y0;
  wire   n2056, n86, n88, n89, n90, n91, n92, n93, n94, n95, n98, n99, n100,
         n101, n103, n104, n107, n108, n109, n110, n112, n113, n115, n116,
         n117, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n136, n152, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n168, n170, n171, n172, n174, n175, n182, n187, n190,
         n191, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n275, n276, n277, n278, n279,
         n280, n281, n283, n284, n285, n291, n296, n297, n298, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n381, n382, n383, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n435, n436, n437, n439, n440, n442, n443, n444, n445,
         n446, n447, n452, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n550, n552, n553, n554, n555,
         n556, n557, n614, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n665, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n688, n690, n691, n695, n696, n697, n701, n702, n703, n704, n709,
         n710, n712, n714, n715, n716, n717, n720, n721, n722, n726, n728,
         n741, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1059, n1060,
         n1062, n1064, n1065, n1066, n1067, n1068, n1069, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1108,
         n1109, n1110, n1111, n1113, n1114, n1115, n1116, n1117, n1118, n1120,
         n1121, n1122, n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135,
         n1136, n1137, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1175, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1238, n1239, n1240, n1241, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1252, n1253, n1254, n1255,
         n1257, n1258, n1259, n1261, n1262, n1263, n1264, n1265, n1266, n1268,
         n1269, n1270, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1280,
         n1281, n1282, n1283, n1284, n1285, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2054, n2055,
         n2057, n2058, n2059, n2060;

  and2 U74 ( .A1(n88), .A2(n89), .Z(n86) );
  or2 U75 ( .A1(n90), .A2(n91), .Z(n89) );
  or2 U76 ( .A1(n92), .A2(n93), .Z(n91) );
  or2 U77 ( .A1(n94), .A2(n95), .Z(n93) );
  and2 U78 ( .A1(q), .A2(n1316), .Z(n95) );
  and2 U79 ( .A1(n2045), .A2(u), .Z(n94) );
  or2 U80 ( .A1(n98), .A2(n99), .Z(n92) );
  and2 U81 ( .A1(n100), .A2(n101), .Z(n99) );
  or2 U82 ( .A1(r), .A2(n2042), .Z(n101) );
  and2 U83 ( .A1(n103), .A2(n104), .Z(n100) );
  or2 U84 ( .A1(s), .A2(n2058), .Z(n103) );
  and2 U85 ( .A1(n2043), .A2(g), .Z(n98) );
  or2 U86 ( .A1(n107), .A2(n108), .Z(n90) );
  or2 U87 ( .A1(n109), .A2(n110), .Z(n108) );
  inv1 U89 ( .I(n112), .ZN(n109) );
  or2 U90 ( .A1(d), .A2(n113), .Z(n107) );
  and2 U91 ( .A1(t), .A2(n2039), .Z(n113) );
  or2 U92 ( .A1(n115), .A2(n116), .Z(n88) );
  or2 U96 ( .A1(n121), .A2(n122), .Z(n117) );
  and2 U97 ( .A1(n2039), .A2(n), .Z(n122) );
  and2 U98 ( .A1(n123), .A2(n124), .Z(n121) );
  or2 U99 ( .A1(m0), .A2(n2058), .Z(n124) );
  and2 U100 ( .A1(n125), .A2(n104), .Z(n123) );
  or2 U101 ( .A1(n0), .A2(n2042), .Z(n125) );
  or2 U102 ( .A1(n126), .A2(n127), .Z(n115) );
  or2 U103 ( .A1(n128), .A2(n129), .Z(n127) );
  or2 U105 ( .A1(n130), .A2(n131), .Z(n126) );
  and2 U106 ( .A1(n2045), .A2(m), .Z(n130) );
  or2 U123 ( .A1(n158), .A2(n159), .Z(n157) );
  or2 U124 ( .A1(n160), .A2(n161), .Z(n159) );
  and2 U125 ( .A1(n162), .A2(n163), .Z(n161) );
  and2 U126 ( .A1(n164), .A2(n165), .Z(n163) );
  inv1 U130 ( .I(n171), .ZN(n164) );
  or2 U131 ( .A1(n172), .A2(n2036), .Z(n171) );
  and2 U132 ( .A1(n174), .A2(n175), .Z(n162) );
  and2 U142 ( .A1(n193), .A2(n194), .Z(n160) );
  and2 U143 ( .A1(n195), .A2(n196), .Z(n194) );
  and2 U144 ( .A1(n197), .A2(n198), .Z(n196) );
  or2 U145 ( .A1(n187), .A2(n199), .Z(n198) );
  or2 U146 ( .A1(n191), .A2(n200), .Z(n197) );
  inv1 U147 ( .I(o), .ZN(n200) );
  and2 U148 ( .A1(n201), .A2(n202), .Z(n195) );
  or2 U149 ( .A1(n203), .A2(n2054), .Z(n202) );
  and2 U151 ( .A1(n207), .A2(n208), .Z(n193) );
  and2 U152 ( .A1(n209), .A2(n210), .Z(n208) );
  or2 U153 ( .A1(n211), .A2(n212), .Z(n210) );
  or2 U154 ( .A1(n2040), .A2(n213), .Z(n212) );
  and2 U155 ( .A1(n2057), .A2(n214), .Z(n213) );
  and2 U156 ( .A1(n182), .A2(n215), .Z(n211) );
  or2 U157 ( .A1(n170), .A2(n216), .Z(n209) );
  and2 U158 ( .A1(n217), .A2(n218), .Z(n207) );
  or2 U159 ( .A1(n219), .A2(n168), .Z(n218) );
  inv1 U160 ( .I(n220), .ZN(n217) );
  and2 U161 ( .A1(n221), .A2(n220), .Z(n158) );
  or2 U162 ( .A1(d), .A2(e), .Z(n220) );
  or2 U213 ( .A1(n276), .A2(n277), .Z(n275) );
  and2 U214 ( .A1(n278), .A2(n279), .Z(n277) );
  and2 U215 ( .A1(n280), .A2(n281), .Z(n279) );
  inv1 U218 ( .I(n284), .ZN(n280) );
  or2 U219 ( .A1(n285), .A2(n2037), .Z(n284) );
  and2 U225 ( .A1(n182), .A2(n190), .Z(n291) );
  inv1 U226 ( .I(m0), .ZN(n190) );
  and2 U231 ( .A1(n296), .A2(n297), .Z(n276) );
  inv1 U235 ( .I(s), .ZN(n216) );
  and2 U236 ( .A1(n301), .A2(n302), .Z(n298) );
  or2 U237 ( .A1(n2051), .A2(n168), .Z(n302) );
  or2 U238 ( .A1(n219), .A2(n2054), .Z(n301) );
  inv1 U240 ( .I(v), .ZN(n219) );
  and2 U241 ( .A1(n303), .A2(n304), .Z(n296) );
  and2 U242 ( .A1(n305), .A2(n306), .Z(n304) );
  inv1 U244 ( .I(u), .ZN(n203) );
  or2 U245 ( .A1(n307), .A2(n308), .Z(n305) );
  or2 U246 ( .A1(n2040), .A2(n309), .Z(n308) );
  and2 U247 ( .A1(n2057), .A2(n199), .Z(n309) );
  inv1 U248 ( .I(r), .ZN(n199) );
  and2 U250 ( .A1(n182), .A2(n214), .Z(n307) );
  inv1 U251 ( .I(q), .ZN(n214) );
  and2 U252 ( .A1(n310), .A2(n311), .Z(n303) );
  or2 U253 ( .A1(n206), .A2(n170), .Z(n311) );
  inv1 U254 ( .I(t), .ZN(n206) );
  or2 U255 ( .A1(n191), .A2(n215), .Z(n310) );
  inv1 U256 ( .I(p), .ZN(n215) );
  and2 U284 ( .A1(n343), .A2(n344), .Z(n342) );
  or2 U285 ( .A1(n345), .A2(n346), .Z(n344) );
  or2 U286 ( .A1(n347), .A2(n348), .Z(n346) );
  or2 U287 ( .A1(n349), .A2(n350), .Z(n348) );
  and2 U288 ( .A1(t), .A2(n1316), .Z(n350) );
  and2 U289 ( .A1(n2045), .A2(h), .Z(n349) );
  or2 U290 ( .A1(n351), .A2(n352), .Z(n347) );
  and2 U291 ( .A1(n353), .A2(n354), .Z(n352) );
  or2 U292 ( .A1(u), .A2(n2042), .Z(n354) );
  and2 U293 ( .A1(n355), .A2(n104), .Z(n353) );
  or2 U294 ( .A1(v), .A2(n2058), .Z(n355) );
  or2 U296 ( .A1(n356), .A2(n357), .Z(n345) );
  or2 U297 ( .A1(n285), .A2(n358), .Z(n357) );
  and2 U298 ( .A1(n2039), .A2(g), .Z(n358) );
  and2 U299 ( .A1(j), .A2(n2043), .Z(n285) );
  or2 U300 ( .A1(d), .A2(n359), .Z(n356) );
  or2 U301 ( .A1(n360), .A2(n361), .Z(n343) );
  or2 U305 ( .A1(n365), .A2(n366), .Z(n362) );
  and2 U306 ( .A1(n2039), .A2(o0), .Z(n366) );
  and2 U307 ( .A1(n367), .A2(n368), .Z(n365) );
  or2 U308 ( .A1(p0), .A2(n2058), .Z(n368) );
  and2 U309 ( .A1(n369), .A2(n104), .Z(n367) );
  or2 U310 ( .A1(q0), .A2(n2042), .Z(n369) );
  or2 U311 ( .A1(n370), .A2(n371), .Z(n360) );
  or2 U312 ( .A1(n372), .A2(n373), .Z(n371) );
  and2 U314 ( .A1(n2043), .A2(n), .Z(n372) );
  or2 U315 ( .A1(n374), .A2(n375), .Z(n370) );
  and2 U316 ( .A1(n2045), .A2(n0), .Z(n374) );
  and2 U318 ( .A1(n378), .A2(n379), .Z(n376) );
  inv1 U320 ( .I(n381), .ZN(n378) );
  or2 U321 ( .A1(n382), .A2(n152), .Z(n381) );
  and2 U337 ( .A1(n402), .A2(n403), .Z(n401) );
  or2 U338 ( .A1(n404), .A2(n405), .Z(n403) );
  or2 U339 ( .A1(n406), .A2(n407), .Z(n405) );
  or2 U340 ( .A1(n408), .A2(n409), .Z(n407) );
  and2 U341 ( .A1(n1316), .A2(u), .Z(n409) );
  and2 U342 ( .A1(n2045), .A2(i), .Z(n408) );
  or2 U343 ( .A1(n410), .A2(n411), .Z(n406) );
  and2 U344 ( .A1(n412), .A2(n413), .Z(n411) );
  or2 U345 ( .A1(g), .A2(n2058), .Z(n413) );
  and2 U346 ( .A1(n414), .A2(n104), .Z(n412) );
  or2 U347 ( .A1(v), .A2(n2042), .Z(n414) );
  and2 U348 ( .A1(n2039), .A2(h), .Z(n410) );
  or2 U349 ( .A1(n415), .A2(n416), .Z(n404) );
  or2 U350 ( .A1(n2036), .A2(n417), .Z(n416) );
  or2 U352 ( .A1(d), .A2(n129), .Z(n415) );
  and2 U353 ( .A1(k), .A2(n2043), .Z(n129) );
  or2 U354 ( .A1(n418), .A2(n419), .Z(n402) );
  or2 U358 ( .A1(n423), .A2(n424), .Z(n420) );
  and2 U359 ( .A1(p0), .A2(n2039), .Z(n424) );
  and2 U360 ( .A1(n425), .A2(n426), .Z(n423) );
  or2 U361 ( .A1(q0), .A2(n2058), .Z(n426) );
  and2 U362 ( .A1(n427), .A2(n104), .Z(n425) );
  or2 U363 ( .A1(r0), .A2(n2042), .Z(n427) );
  or2 U364 ( .A1(n428), .A2(n429), .Z(n418) );
  or2 U365 ( .A1(n430), .A2(n431), .Z(n429) );
  and2 U366 ( .A1(n2043), .A2(m0), .Z(n431) );
  or2 U368 ( .A1(n432), .A2(n433), .Z(n428) );
  and2 U369 ( .A1(n2044), .A2(n), .Z(n433) );
  and2 U370 ( .A1(n2045), .A2(o0), .Z(n432) );
  and2 U372 ( .A1(n436), .A2(n437), .Z(n435) );
  and2 U374 ( .A1(n439), .A2(n440), .Z(n436) );
  or2 U376 ( .A1(n443), .A2(n444), .Z(n442) );
  and2 U377 ( .A1(n445), .A2(f), .Z(n444) );
  and2 U378 ( .A1(n446), .A2(n447), .Z(n443) );
  or2 U383 ( .A1(n152), .A2(n452), .Z(n439) );
  and2 U392 ( .A1(n462), .A2(n463), .Z(n461) );
  or2 U393 ( .A1(n464), .A2(n465), .Z(n463) );
  or2 U394 ( .A1(n466), .A2(n467), .Z(n465) );
  or2 U395 ( .A1(n468), .A2(n469), .Z(n467) );
  and2 U396 ( .A1(s), .A2(n1316), .Z(n469) );
  and2 U397 ( .A1(n2039), .A2(v), .Z(n468) );
  or2 U398 ( .A1(n470), .A2(n471), .Z(n466) );
  and2 U399 ( .A1(n472), .A2(n473), .Z(n471) );
  or2 U400 ( .A1(t), .A2(n2042), .Z(n473) );
  and2 U401 ( .A1(n474), .A2(n104), .Z(n472) );
  or2 U402 ( .A1(u), .A2(n2058), .Z(n474) );
  or2 U404 ( .A1(n475), .A2(n476), .Z(n464) );
  or2 U405 ( .A1(n172), .A2(n477), .Z(n476) );
  and2 U406 ( .A1(n2045), .A2(g), .Z(n477) );
  and2 U407 ( .A1(i), .A2(n2043), .Z(n172) );
  or2 U408 ( .A1(d), .A2(n131), .Z(n475) );
  and2 U409 ( .A1(j), .A2(n2044), .Z(n131) );
  or2 U410 ( .A1(n478), .A2(n479), .Z(n462) );
  or2 U414 ( .A1(n483), .A2(n484), .Z(n480) );
  and2 U415 ( .A1(n2039), .A2(n0), .Z(n484) );
  and2 U416 ( .A1(n485), .A2(n486), .Z(n483) );
  or2 U417 ( .A1(o0), .A2(n2058), .Z(n486) );
  and2 U418 ( .A1(n487), .A2(n104), .Z(n485) );
  or2 U419 ( .A1(p0), .A2(n2042), .Z(n487) );
  or2 U420 ( .A1(n488), .A2(n489), .Z(n478) );
  or2 U421 ( .A1(n490), .A2(n491), .Z(n489) );
  and2 U422 ( .A1(n2043), .A2(m), .Z(n491) );
  or2 U424 ( .A1(n492), .A2(n417), .Z(n488) );
  and2 U425 ( .A1(l), .A2(n2044), .Z(n417) );
  and2 U426 ( .A1(n2045), .A2(m0), .Z(n492) );
  and2 U428 ( .A1(n494), .A2(n495), .Z(n493) );
  inv1 U430 ( .I(n496), .ZN(n494) );
  or2 U431 ( .A1(n497), .A2(n152), .Z(n496) );
  or2 U475 ( .A1(n552), .A2(n553), .Z(n550) );
  and2 U476 ( .A1(i), .A2(n2051), .Z(n553) );
  and2 U477 ( .A1(j), .A2(n554), .Z(n552) );
  or2 U478 ( .A1(n555), .A2(n556), .Z(n554) );
  and2 U479 ( .A1(i), .A2(n2050), .Z(n556) );
  and2 U480 ( .A1(n557), .A2(g), .Z(n555) );
  and2 U481 ( .A1(h), .A2(n2049), .Z(n557) );
  and2 U536 ( .A1(n617), .A2(n618), .Z(n616) );
  or2 U537 ( .A1(n619), .A2(n620), .Z(n618) );
  or2 U538 ( .A1(n621), .A2(n622), .Z(n620) );
  or2 U539 ( .A1(n623), .A2(n624), .Z(n622) );
  and2 U540 ( .A1(n1316), .A2(r), .Z(n624) );
  and2 U541 ( .A1(n2045), .A2(v), .Z(n623) );
  or2 U542 ( .A1(n625), .A2(n626), .Z(n621) );
  and2 U543 ( .A1(n627), .A2(n628), .Z(n626) );
  or2 U544 ( .A1(s), .A2(n2042), .Z(n628) );
  and2 U545 ( .A1(n629), .A2(n104), .Z(n627) );
  or2 U546 ( .A1(t), .A2(n2058), .Z(n629) );
  or2 U548 ( .A1(n630), .A2(n631), .Z(n619) );
  or2 U549 ( .A1(n632), .A2(n633), .Z(n631) );
  and2 U550 ( .A1(n2043), .A2(h), .Z(n633) );
  inv1 U551 ( .I(n283), .ZN(n632) );
  or2 U553 ( .A1(d), .A2(n634), .Z(n630) );
  and2 U554 ( .A1(n2039), .A2(u), .Z(n634) );
  or2 U555 ( .A1(n635), .A2(n636), .Z(n617) );
  or2 U559 ( .A1(n640), .A2(n641), .Z(n637) );
  and2 U560 ( .A1(n2045), .A2(n), .Z(n641) );
  and2 U561 ( .A1(n642), .A2(n643), .Z(n640) );
  or2 U562 ( .A1(n0), .A2(n2058), .Z(n643) );
  and2 U563 ( .A1(n644), .A2(n104), .Z(n642) );
  or2 U564 ( .A1(o0), .A2(n2042), .Z(n644) );
  or2 U565 ( .A1(n645), .A2(n646), .Z(n635) );
  or2 U566 ( .A1(n647), .A2(n648), .Z(n646) );
  or2 U568 ( .A1(n649), .A2(n359), .Z(n645) );
  and2 U569 ( .A1(k), .A2(n2044), .Z(n359) );
  and2 U570 ( .A1(n2039), .A2(m0), .Z(n649) );
  or2 U571 ( .A1(j), .A2(n132), .Z(n614) );
  and2 U589 ( .A1(n668), .A2(n669), .Z(n667) );
  or2 U590 ( .A1(n670), .A2(n671), .Z(n669) );
  or2 U591 ( .A1(n672), .A2(n673), .Z(n671) );
  or2 U592 ( .A1(n674), .A2(n675), .Z(n673) );
  and2 U593 ( .A1(n1316), .A2(v), .Z(n675) );
  and2 U594 ( .A1(n2045), .A2(j), .Z(n674) );
  or2 U595 ( .A1(n676), .A2(n677), .Z(n672) );
  and2 U596 ( .A1(n678), .A2(n679), .Z(n677) );
  or2 U597 ( .A1(g), .A2(n2042), .Z(n679) );
  and2 U598 ( .A1(n680), .A2(n104), .Z(n678) );
  or2 U599 ( .A1(h), .A2(n2058), .Z(n680) );
  and2 U600 ( .A1(n2039), .A2(i), .Z(n676) );
  or2 U601 ( .A1(n681), .A2(n682), .Z(n670) );
  or2 U602 ( .A1(n2037), .A2(n375), .Z(n682) );
  and2 U603 ( .A1(m), .A2(n2044), .Z(n375) );
  or2 U605 ( .A1(d), .A2(n648), .Z(n681) );
  and2 U606 ( .A1(l), .A2(n2043), .Z(n648) );
  or2 U607 ( .A1(n683), .A2(n684), .Z(n668) );
  or2 U613 ( .A1(n690), .A2(n691), .Z(n685) );
  and2 U614 ( .A1(q0), .A2(n2039), .Z(n691) );
  and2 U618 ( .A1(n695), .A2(n696), .Z(n690) );
  or2 U619 ( .A1(r0), .A2(n2058), .Z(n696) );
  and2 U620 ( .A1(n697), .A2(n104), .Z(n695) );
  or2 U625 ( .A1(s0), .A2(n2042), .Z(n697) );
  or2 U628 ( .A1(n701), .A2(n702), .Z(n683) );
  or2 U629 ( .A1(n703), .A2(n704), .Z(n702) );
  and2 U630 ( .A1(n2043), .A2(n0), .Z(n704) );
  or2 U638 ( .A1(n709), .A2(n710), .Z(n701) );
  and2 U639 ( .A1(n2044), .A2(m0), .Z(n710) );
  and2 U644 ( .A1(p0), .A2(n2045), .Z(n709) );
  or2 U647 ( .A1(z), .A2(y), .Z(n688) );
  or2 U649 ( .A1(n712), .A2(n377), .Z(n665) );
  and2 U653 ( .A1(c), .A2(n715), .Z(n714) );
  and2 U654 ( .A1(n716), .A2(n717), .Z(n712) );
  and2 U659 ( .A1(n720), .A2(n721), .Z(n716) );
  or2 U660 ( .A1(n152), .A2(n722), .Z(n721) );
  or2 U666 ( .A1(f), .A2(n2047), .Z(n726) );
  inv1 U672 ( .I(n136), .ZN(n152) );
  or2 U673 ( .A1(b), .A2(d), .Z(n136) );
  and2 U686 ( .A1(n2047), .A2(n2046), .Z(n741) );
  and2 U1051 ( .A1(n1051), .A2(n1052), .Z(c1) );
  inv1 U1052 ( .I(n1053), .ZN(n1052) );
  and2 U1053 ( .A1(n728), .A2(n383), .Z(n1053) );
  or2 U1054 ( .A1(n383), .A2(n728), .Z(n1051) );
  and2 U1055 ( .A1(n1054), .A2(n1055), .Z(n728) );
  and2 U1057 ( .A1(n1057), .A2(n2048), .Z(n1056) );
  or2 U1058 ( .A1(n2048), .A2(n1057), .Z(n1054) );
  or2 U1059 ( .A1(n1059), .A2(n1060), .Z(n1057) );
  and2 U1060 ( .A1(g), .A2(n2050), .Z(n1060) );
  and2 U1061 ( .A1(h), .A2(n2051), .Z(n1059) );
  and2 U1065 ( .A1(j), .A2(n2049), .Z(n1062) );
  or2 U1066 ( .A1(n1064), .A2(n1065), .Z(n383) );
  and2 U1067 ( .A1(n1066), .A2(n1067), .Z(n1065) );
  and2 U1069 ( .A1(n1068), .A2(n1069), .Z(n1064) );
  and2 U1077 ( .A1(n1074), .A2(n1075), .Z(b1) );
  inv1 U1078 ( .I(n1076), .ZN(n1075) );
  and2 U1079 ( .A1(n445), .A2(n498), .Z(n1076) );
  or2 U1080 ( .A1(n498), .A2(n445), .Z(n1074) );
  and2 U1081 ( .A1(n1077), .A2(n1078), .Z(n445) );
  inv1 U1082 ( .I(n1079), .ZN(n1078) );
  and2 U1083 ( .A1(n1080), .A2(n1081), .Z(n1079) );
  or2 U1084 ( .A1(n1081), .A2(n1080), .Z(n1077) );
  or2 U1085 ( .A1(n1082), .A2(n1083), .Z(n1080) );
  and2 U1086 ( .A1(d0), .A2(n1084), .Z(n1083) );
  and2 U1087 ( .A1(e0), .A2(n1085), .Z(n1082) );
  inv1 U1088 ( .I(n1086), .ZN(n1081) );
  or2 U1089 ( .A1(n1087), .A2(n1088), .Z(n1086) );
  and2 U1090 ( .A1(f0), .A2(n1089), .Z(n1088) );
  and2 U1091 ( .A1(g0), .A2(n1090), .Z(n1087) );
  or2 U1092 ( .A1(n1091), .A2(n1092), .Z(n498) );
  and2 U1093 ( .A1(n1093), .A2(n1094), .Z(n1092) );
  inv1 U1094 ( .I(n1095), .ZN(n1094) );
  and2 U1095 ( .A1(n1095), .A2(n1096), .Z(n1091) );
  inv1 U1096 ( .I(n1093), .ZN(n1096) );
  or2 U1097 ( .A1(n1097), .A2(n1098), .Z(n1093) );
  and2 U1098 ( .A1(h0), .A2(n1099), .Z(n1098) );
  and2 U1099 ( .A1(i0), .A2(n1100), .Z(n1097) );
  or2 U1100 ( .A1(n1101), .A2(n1102), .Z(n1095) );
  and2 U1101 ( .A1(j0), .A2(n1103), .Z(n1102) );
  and2 U1102 ( .A1(k0), .A2(n1104), .Z(n1101) );
  and2 U1103 ( .A1(n1105), .A2(n2055), .Z(a1) );
  and2 U1108 ( .A1(n1108), .A2(n1109), .Z(n1105) );
  or2 U1109 ( .A1(n1110), .A2(n1111), .Z(n1109) );
  and2 U1112 ( .A1(n1113), .A2(n1114), .Z(n1110) );
  and2 U1113 ( .A1(n1115), .A2(n1116), .Z(n1114) );
  and2 U1114 ( .A1(n1117), .A2(n1118), .Z(n1116) );
  or2 U1115 ( .A1(n2051), .A2(n1085), .Z(n1118) );
  inv1 U1116 ( .I(d0), .ZN(n1085) );
  or2 U1118 ( .A1(n2050), .A2(n1084), .Z(n1117) );
  inv1 U1119 ( .I(e0), .ZN(n1084) );
  or2 U1122 ( .A1(n1090), .A2(n2049), .Z(n1120) );
  inv1 U1124 ( .I(f0), .ZN(n1090) );
  inv1 U1126 ( .I(g0), .ZN(n1089) );
  and2 U1128 ( .A1(n1121), .A2(n1122), .Z(n1113) );
  inv1 U1138 ( .I(k0), .ZN(n1103) );
  or2 U1140 ( .A1(n1100), .A2(n1127), .Z(n1108) );
  and2 U1146 ( .A1(n1099), .A2(n1104), .Z(n1128) );
  inv1 U1147 ( .I(j0), .ZN(n1104) );
  inv1 U1148 ( .I(i0), .ZN(n1099) );
  inv1 U1149 ( .I(h0), .ZN(n1100) );
  or2 U1154 ( .A1(e), .A2(a), .Z(n1133) );
  or2 U1158 ( .A1(n1212), .A2(n1634), .Z(n1136) );
  or2 U1159 ( .A1(n1233), .A2(n1137), .Z(n1244) );
  or2 U1160 ( .A1(n1129), .A2(n1979), .Z(n1137) );
  inv1 U1163 ( .I(n1719), .ZN(n1140) );
  and2 U1167 ( .A1(n1152), .A2(n1449), .Z(n1143) );
  or2 U1168 ( .A1(d), .A2(w0), .Z(n1144) );
  and2 U1169 ( .A1(n1671), .A2(n1670), .Z(n1145) );
  inv1 U1170 ( .I(n1145), .ZN(n1682) );
  inv1 U1172 ( .I(n1146), .ZN(n2022) );
  and2 U1179 ( .A1(n1152), .A2(n1449), .Z(n1151) );
  inv1 U1180 ( .I(n1471), .ZN(n1152) );
  and2 U1181 ( .A1(n1201), .A2(n1504), .Z(n1153) );
  and2 U1182 ( .A1(n1195), .A2(n1155), .Z(n1154) );
  inv1 U1183 ( .I(n1223), .ZN(n1155) );
  and2 U1184 ( .A1(n1181), .A2(n1394), .Z(n1156) );
  and2 U1187 ( .A1(i0), .A2(n1159), .Z(n1158) );
  inv1 U1188 ( .I(n1456), .ZN(n1159) );
  inv1 U1189 ( .I(a), .ZN(n1160) );
  and2 U1192 ( .A1(n1445), .A2(n1446), .Z(n1163) );
  or2 U1193 ( .A1(n1163), .A2(n1164), .Z(n1449) );
  or2 U1194 ( .A1(n1448), .A2(n1447), .Z(n1164) );
  inv1 U1195 ( .I(n1383), .ZN(n1165) );
  and2 U1196 ( .A1(c), .A2(d), .Z(n1166) );
  or2 U1197 ( .A1(n1872), .A2(n1169), .Z(n1167) );
  or2 U1200 ( .A1(n1873), .A2(n1905), .Z(n1169) );
  and2 U1201 ( .A1(n1863), .A2(n1898), .Z(n1170) );
  and2 U1203 ( .A1(e), .A2(d), .Z(n1172) );
  or2 U1209 ( .A1(n1172), .A2(n1179), .Z(n1178) );
  or2 U1212 ( .A1(n1203), .A2(b), .Z(n1181) );
  and2 U1213 ( .A1(n1762), .A2(n1763), .Z(n1182) );
  or2 U1215 ( .A1(n1898), .A2(n1765), .Z(n1183) );
  or2 U1216 ( .A1(n1419), .A2(n1418), .Z(n1184) );
  or2 U1223 ( .A1(n1639), .A2(n1191), .Z(n1189) );
  and2 U1224 ( .A1(n1189), .A2(n1190), .Z(n1640) );
  or2 U1225 ( .A1(n1757), .A2(n1735), .Z(n1190) );
  or2 U1226 ( .A1(n1252), .A2(n1757), .Z(n1191) );
  and2 U1227 ( .A1(b), .A2(a), .Z(n1192) );
  and2 U1228 ( .A1(n1614), .A2(n1613), .Z(n1193) );
  inv1 U1229 ( .I(n1180), .ZN(n1282) );
  inv1 U1230 ( .I(n1431), .ZN(n1194) );
  inv1 U1232 ( .I(n1224), .ZN(n1196) );
  or2 U1233 ( .A1(n1501), .A2(n1499), .Z(n1197) );
  or2 U1234 ( .A1(n1642), .A2(n1641), .Z(n1198) );
  or2 U1235 ( .A1(n1193), .A2(n1248), .Z(n1199) );
  inv1 U1237 ( .I(n1200), .ZN(n1466) );
  or2 U1238 ( .A1(n1210), .A2(n1211), .Z(n1201) );
  and2 U1240 ( .A1(c), .A2(d), .Z(n1203) );
  and2 U1245 ( .A1(b), .A2(a), .Z(n1207) );
  or2 U1246 ( .A1(n1561), .A2(n1562), .Z(n1208) );
  inv1 U1248 ( .I(n1489), .ZN(n1210) );
  inv1 U1249 ( .I(n1488), .ZN(n1211) );
  inv1 U1250 ( .I(n1247), .ZN(n1212) );
  and2 U1251 ( .A1(n1524), .A2(g0), .Z(n1213) );
  or2 U1252 ( .A1(n1717), .A2(n1216), .Z(n1214) );
  or2 U1254 ( .A1(n1724), .A2(n1941), .Z(n1215) );
  or2 U1255 ( .A1(n1716), .A2(n1724), .Z(n1216) );
  and2 U1257 ( .A1(n1209), .A2(n1504), .Z(n1218) );
  and2 U1258 ( .A1(u0), .A2(n1713), .Z(n1219) );
  inv1 U1259 ( .I(n2025), .ZN(n1220) );
  and2 U1263 ( .A1(n1225), .A2(n1219), .Z(n1223) );
  and2 U1264 ( .A1(n1711), .A2(u0), .Z(n1224) );
  and2 U1267 ( .A1(n1226), .A2(n1227), .Z(n1883) );
  or2 U1268 ( .A1(n1881), .A2(n1880), .Z(n1227) );
  or2 U1269 ( .A1(n1878), .A2(n1881), .Z(n1228) );
  inv1 U1271 ( .I(n1229), .ZN(n1243) );
  inv1 U1272 ( .I(n1280), .ZN(n1230) );
  inv1 U1273 ( .I(n1254), .ZN(n1231) );
  or2 U1281 ( .A1(n1687), .A2(n1238), .Z(n1239) );
  or2 U1282 ( .A1(n1686), .A2(n1878), .Z(n1238) );
  inv1 U1283 ( .I(n1239), .ZN(n1716) );
  or2 U1284 ( .A1(n1869), .A2(n1154), .Z(n1240) );
  or2 U1287 ( .A1(n1611), .A2(n1610), .Z(n1245) );
  or2 U1288 ( .A1(n1506), .A2(n1153), .Z(n1246) );
  or2 U1289 ( .A1(n1626), .A2(n1248), .Z(n1247) );
  inv1 U1290 ( .I(n1199), .ZN(n1252) );
  inv1 U1291 ( .I(n1625), .ZN(n1248) );
  and2 U1292 ( .A1(n1510), .A2(n1509), .Z(n1249) );
  or2 U1296 ( .A1(n1507), .A2(n1881), .Z(n1253) );
  or2 U1303 ( .A1(n1259), .A2(n1869), .Z(n1870) );
  or2 U1304 ( .A1(n1154), .A2(n1875), .Z(n1259) );
  or2 U1308 ( .A1(n1161), .A2(n1409), .Z(n1262) );
  or2 U1310 ( .A1(n1240), .A2(n1875), .Z(n1264) );
  or2 U1312 ( .A1(n1486), .A2(n1487), .Z(n1266) );
  and2 U1317 ( .A1(b), .A2(a), .Z(n1270) );
  or2 U1322 ( .A1(n1982), .A2(x0), .Z(n1275) );
  inv1 U1324 ( .I(n1265), .ZN(n1278) );
  or2 U1326 ( .A1(n1282), .A2(n1437), .Z(n1280) );
  inv1 U1327 ( .I(n1995), .ZN(n1283) );
  inv1 U1328 ( .I(d), .ZN(n1285) );
  inv1 U1329 ( .I(d), .ZN(n1284) );
  or2 U1332 ( .A1(b), .A2(n1160), .Z(n1775) );
  inv1 U1333 ( .I(c), .ZN(n1695) );
  or2 U1334 ( .A1(n1775), .A2(n1695), .Z(n1302) );
  or2 U1335 ( .A1(n1302), .A2(n1128), .Z(n1127) );
  inv1 U1336 ( .I(m), .ZN(n1493) );
  or2 U1337 ( .A1(n1104), .A2(n1493), .Z(n1288) );
  inv1 U1338 ( .I(n), .ZN(n1444) );
  or2 U1339 ( .A1(n1103), .A2(n1444), .Z(n1287) );
  and2 U1340 ( .A1(n1288), .A2(n1287), .Z(n1121) );
  inv1 U1341 ( .I(k), .ZN(n1421) );
  or2 U1342 ( .A1(n1100), .A2(n1421), .Z(n1290) );
  inv1 U1343 ( .I(l), .ZN(n1395) );
  or2 U1344 ( .A1(n1099), .A2(n1395), .Z(n1289) );
  and2 U1345 ( .A1(n1290), .A2(n1289), .Z(n1122) );
  inv1 U1346 ( .I(i), .ZN(n2049) );
  inv1 U1347 ( .I(h), .ZN(n2050) );
  inv1 U1348 ( .I(g), .ZN(n2051) );
  inv1 U1349 ( .I(j), .ZN(n1547) );
  or2 U1350 ( .A1(n1089), .A2(n1547), .Z(n1291) );
  and2 U1351 ( .A1(n1120), .A2(n1291), .Z(n1115) );
  or2 U1352 ( .A1(n1205), .A2(n1695), .Z(n1292) );
  or2 U1353 ( .A1(n1292), .A2(n1160), .Z(n1728) );
  inv1 U1354 ( .I(n1728), .ZN(n1781) );
  inv1 U1355 ( .I(n1302), .ZN(n1293) );
  or2 U1356 ( .A1(n1781), .A2(n1293), .Z(n1111) );
  or2 U1357 ( .A1(i), .A2(h), .Z(n1515) );
  inv1 U1358 ( .I(n1515), .ZN(n1576) );
  or2 U1359 ( .A1(n1728), .A2(n2051), .Z(n1294) );
  or2 U1360 ( .A1(n1576), .A2(n1294), .Z(n2055) );
  and2 U1361 ( .A1(n), .A2(n1493), .Z(n1296) );
  and2 U1362 ( .A1(n1444), .A2(m), .Z(n1295) );
  or2 U1363 ( .A1(n1296), .A2(n1295), .Z(n1068) );
  and2 U1364 ( .A1(l), .A2(n1421), .Z(n1298) );
  and2 U1365 ( .A1(n1395), .A2(k), .Z(n1297) );
  or2 U1366 ( .A1(n1298), .A2(n1297), .Z(n1066) );
  inv1 U1367 ( .I(n1066), .ZN(n1069) );
  inv1 U1368 ( .I(n1068), .ZN(n1067) );
  and2 U1369 ( .A1(n1547), .A2(i), .Z(n1299) );
  or2 U1370 ( .A1(n1299), .A2(n1062), .Z(n1300) );
  inv1 U1371 ( .I(n1300), .ZN(n2048) );
  inv1 U1372 ( .I(n1056), .ZN(n1055) );
  or2 U1373 ( .A1(n1576), .A2(n2051), .Z(n1301) );
  inv1 U1374 ( .I(n1301), .ZN(n2047) );
  or2 U1375 ( .A1(n1302), .A2(e), .Z(n1905) );
  inv1 U1376 ( .I(n1905), .ZN(n2046) );
  or2 U1377 ( .A1(n1302), .A2(n1285), .Z(n1328) );
  inv1 U1378 ( .I(n1328), .ZN(n1333) );
  or2 U1379 ( .A1(n1333), .A2(n), .Z(n722) );
  or2 U1381 ( .A1(n728), .A2(n1527), .Z(n1303) );
  and2 U1382 ( .A1(n726), .A2(n1303), .Z(n1304) );
  or2 U1383 ( .A1(n1304), .A2(n1328), .Z(n720) );
  or2 U1384 ( .A1(m), .A2(l), .Z(n1324) );
  inv1 U1385 ( .I(n1324), .ZN(n1305) );
  or2 U1386 ( .A1(n1305), .A2(n1421), .Z(z0) );
  inv1 U1387 ( .I(z0), .ZN(n1306) );
  or2 U1388 ( .A1(n1306), .A2(n136), .Z(n717) );
  inv1 U1389 ( .I(w), .ZN(n715) );
  and2 U1390 ( .A1(n152), .A2(n1695), .Z(n1702) );
  or2 U1391 ( .A1(n1205), .A2(n714), .Z(n1937) );
  inv1 U1392 ( .I(n1937), .ZN(n1925) );
  or2 U1393 ( .A1(n1702), .A2(n1925), .Z(n377) );
  inv1 U1394 ( .I(x), .ZN(n1612) );
  or2 U1395 ( .A1(n1695), .A2(n1612), .Z(n1313) );
  or2 U1396 ( .A1(n1313), .A2(n688), .Z(n170) );
  inv1 U1397 ( .I(n170), .ZN(n2045) );
  inv1 U1398 ( .I(z), .ZN(n1628) );
  or2 U1399 ( .A1(n1695), .A2(n1628), .Z(n1307) );
  or2 U1400 ( .A1(n1307), .A2(x), .Z(n1309) );
  or2 U1401 ( .A1(n1309), .A2(y), .Z(n168) );
  inv1 U1402 ( .I(n168), .ZN(n2044) );
  inv1 U1403 ( .I(y), .ZN(n1630) );
  or2 U1404 ( .A1(z), .A2(n1630), .Z(n1310) );
  and2 U1405 ( .A1(c), .A2(n1310), .Z(n1308) );
  inv1 U1406 ( .I(n1313), .ZN(n1312) );
  or2 U1407 ( .A1(n1308), .A2(n1312), .Z(n2054) );
  inv1 U1408 ( .I(n2054), .ZN(n2043) );
  or2 U1409 ( .A1(n1309), .A2(n1630), .Z(n1348) );
  inv1 U1410 ( .I(n1348), .ZN(n1361) );
  and2 U1411 ( .A1(o0), .A2(n1361), .Z(n703) );
  or2 U1412 ( .A1(n1310), .A2(n1313), .Z(n182) );
  and2 U1414 ( .A1(y), .A2(z), .Z(n1311) );
  and2 U1415 ( .A1(n1312), .A2(n1311), .Z(n2041) );
  or2 U1417 ( .A1(n1313), .A2(n1628), .Z(n1314) );
  or2 U1418 ( .A1(n1314), .A2(y), .Z(n187) );
  inv1 U1419 ( .I(n187), .ZN(n2039) );
  or2 U1420 ( .A1(n1695), .A2(n688), .Z(n1315) );
  or2 U1421 ( .A1(n1315), .A2(x), .Z(n191) );
  inv1 U1422 ( .I(n191), .ZN(n1316) );
  and2 U1423 ( .A1(n1316), .A2(t0), .Z(n1317) );
  or2 U1424 ( .A1(n1285), .A2(n1317), .Z(n1318) );
  or2 U1425 ( .A1(n685), .A2(n1318), .Z(n684) );
  or2 U1426 ( .A1(n1348), .A2(n1421), .Z(n1319) );
  inv1 U1427 ( .I(n1319), .ZN(n2037) );
  or2 U1429 ( .A1(n1925), .A2(n152), .Z(n132) );
  and2 U1430 ( .A1(m), .A2(n1361), .Z(n647) );
  and2 U1431 ( .A1(n1316), .A2(p0), .Z(n1320) );
  or2 U1432 ( .A1(n1285), .A2(n1320), .Z(n1321) );
  or2 U1433 ( .A1(n637), .A2(n1321), .Z(n636) );
  or2 U1434 ( .A1(n168), .A2(n2049), .Z(n283) );
  and2 U1435 ( .A1(g), .A2(n1361), .Z(n625) );
  and2 U1436 ( .A1(n498), .A2(n1333), .Z(n497) );
  or2 U1437 ( .A1(n1333), .A2(k), .Z(n495) );
  and2 U1438 ( .A1(n), .A2(n1361), .Z(n490) );
  and2 U1439 ( .A1(n1316), .A2(q0), .Z(n1322) );
  or2 U1440 ( .A1(n1285), .A2(n1322), .Z(n1323) );
  or2 U1441 ( .A1(n480), .A2(n1323), .Z(n479) );
  and2 U1442 ( .A1(h), .A2(n1361), .Z(n470) );
  or2 U1443 ( .A1(n1333), .A2(m), .Z(n452) );
  or2 U1444 ( .A1(n1324), .A2(k), .Z(n1426) );
  or2 U1445 ( .A1(n1426), .A2(n), .Z(n1688) );
  or2 U1446 ( .A1(n1688), .A2(n2050), .Z(n1325) );
  inv1 U1447 ( .I(n1325), .ZN(n446) );
  and2 U1448 ( .A1(n1527), .A2(n2051), .Z(n1327) );
  or2 U1449 ( .A1(n2049), .A2(n1547), .Z(n1326) );
  and2 U1450 ( .A1(n1327), .A2(n1326), .Z(n447) );
  or2 U1451 ( .A1(n1328), .A2(n442), .Z(n440) );
  and2 U1452 ( .A1(n152), .A2(n1688), .Z(n1329) );
  inv1 U1453 ( .I(n1329), .ZN(n437) );
  and2 U1454 ( .A1(n0), .A2(n1361), .Z(n430) );
  and2 U1455 ( .A1(n1316), .A2(s0), .Z(n1330) );
  or2 U1456 ( .A1(n1285), .A2(n1330), .Z(n1331) );
  or2 U1457 ( .A1(n420), .A2(n1331), .Z(n419) );
  or2 U1458 ( .A1(n1348), .A2(n1547), .Z(n1332) );
  inv1 U1459 ( .I(n1332), .ZN(n2036) );
  and2 U1460 ( .A1(n383), .A2(n1333), .Z(n382) );
  or2 U1461 ( .A1(n1333), .A2(l), .Z(n379) );
  and2 U1462 ( .A1(m0), .A2(n1361), .Z(n373) );
  and2 U1463 ( .A1(n1316), .A2(r0), .Z(n1334) );
  or2 U1464 ( .A1(n1285), .A2(n1334), .Z(n1335) );
  or2 U1465 ( .A1(n362), .A2(n1335), .Z(n361) );
  and2 U1466 ( .A1(i), .A2(n1361), .Z(n351) );
  inv1 U1467 ( .I(n104), .ZN(n2040) );
  or2 U1468 ( .A1(n1348), .A2(n203), .Z(n306) );
  and2 U1469 ( .A1(n298), .A2(n1285), .Z(n1337) );
  or2 U1470 ( .A1(n187), .A2(n216), .Z(n1336) );
  and2 U1471 ( .A1(n1337), .A2(n1336), .Z(n297) );
  or2 U1472 ( .A1(n170), .A2(n1395), .Z(n1338) );
  and2 U1473 ( .A1(n283), .A2(n1338), .Z(n281) );
  or2 U1474 ( .A1(n2058), .A2(n), .Z(n1339) );
  inv1 U1475 ( .I(n1339), .ZN(n1340) );
  or2 U1476 ( .A1(n1340), .A2(n2040), .Z(n1341) );
  or2 U1477 ( .A1(n1341), .A2(n291), .Z(n1342) );
  and2 U1478 ( .A1(d), .A2(n1342), .Z(n1347) );
  inv1 U1479 ( .I(n0), .ZN(n1343) );
  or2 U1480 ( .A1(n191), .A2(n1343), .Z(n1345) );
  or2 U1481 ( .A1(n187), .A2(n1493), .Z(n1344) );
  and2 U1482 ( .A1(n1345), .A2(n1344), .Z(n1346) );
  and2 U1483 ( .A1(n1347), .A2(n1346), .Z(n278) );
  or2 U1484 ( .A1(e), .A2(n1285), .Z(n1349) );
  and2 U1485 ( .A1(n2051), .A2(n1349), .Z(n221) );
  or2 U1486 ( .A1(n1348), .A2(n206), .Z(n201) );
  inv1 U1487 ( .I(n1349), .ZN(n1351) );
  or2 U1488 ( .A1(n191), .A2(n190), .Z(n1350) );
  and2 U1489 ( .A1(n1351), .A2(n1350), .Z(n174) );
  or2 U1490 ( .A1(n2058), .A2(m), .Z(n1352) );
  inv1 U1491 ( .I(n1352), .ZN(n1355) );
  and2 U1492 ( .A1(n1444), .A2(n182), .Z(n1353) );
  or2 U1493 ( .A1(n1353), .A2(n2040), .Z(n1354) );
  or2 U1494 ( .A1(n1355), .A2(n1354), .Z(n1357) );
  or2 U1495 ( .A1(n187), .A2(n1395), .Z(n1356) );
  and2 U1496 ( .A1(n1357), .A2(n1356), .Z(n175) );
  or2 U1497 ( .A1(n168), .A2(n2050), .Z(n112) );
  or2 U1498 ( .A1(n170), .A2(n1421), .Z(n1358) );
  and2 U1499 ( .A1(n112), .A2(n1358), .Z(n165) );
  and2 U1500 ( .A1(l), .A2(n1361), .Z(n128) );
  and2 U1501 ( .A1(n1316), .A2(o0), .Z(n1359) );
  or2 U1502 ( .A1(n1285), .A2(n1359), .Z(n1360) );
  or2 U1503 ( .A1(n117), .A2(n1360), .Z(n116) );
  and2 U1504 ( .A1(v), .A2(n1361), .Z(n110) );
  or2 U1505 ( .A1(n1515), .A2(g), .Z(n1362) );
  or2 U1506 ( .A1(n1362), .A2(j), .Z(n1363) );
  inv1 U1507 ( .I(n1363), .ZN(y0) );
  or2 U1508 ( .A1(d), .A2(w0), .Z(n1456) );
  or2 U1509 ( .A1(n1144), .A2(n1177), .Z(n1364) );
  inv1 U1512 ( .I(l0), .ZN(n1528) );
  or2 U1514 ( .A1(n1528), .A2(n1365), .Z(n1366) );
  or2 U1515 ( .A1(n1366), .A2(e), .Z(n1367) );
  inv1 U1516 ( .I(n1367), .ZN(n1480) );
  and2 U1520 ( .A1(m0), .A2(n1601), .Z(n1377) );
  inv1 U1521 ( .I(w0), .ZN(n1370) );
  and2 U1524 ( .A1(n1171), .A2(h0), .Z(n1375) );
  or2 U1525 ( .A1(e), .A2(a), .Z(n1372) );
  and2 U1527 ( .A1(n1482), .A2(i0), .Z(n1373) );
  and2 U1528 ( .A1(n1281), .A2(n1373), .Z(n1374) );
  or2 U1531 ( .A1(n1378), .A2(n1379), .Z(n1680) );
  or2 U1532 ( .A1(n1254), .A2(n1612), .Z(n1381) );
  inv1 U1533 ( .I(n1680), .ZN(n1673) );
  or2 U1534 ( .A1(n1673), .A2(n715), .Z(n1380) );
  or2 U1536 ( .A1(n1186), .A2(l), .Z(n1389) );
  or2 U1537 ( .A1(n1166), .A2(b), .Z(n1383) );
  and2 U1538 ( .A1(a), .A2(n1383), .Z(n1386) );
  and2 U1539 ( .A1(d), .A2(n2059), .Z(n1384) );
  or2 U1542 ( .A1(n1263), .A2(n1395), .Z(n1388) );
  and2 U1543 ( .A1(n1389), .A2(n1388), .Z(n1392) );
  or2 U1544 ( .A1(c), .A2(n1285), .Z(n1438) );
  inv1 U1547 ( .I(n1390), .ZN(n1619) );
  and2 U1548 ( .A1(m), .A2(n1619), .Z(n1391) );
  or2 U1549 ( .A1(n1392), .A2(n1391), .Z(n1402) );
  or2 U1550 ( .A1(c), .A2(d), .Z(n1440) );
  and2 U1553 ( .A1(j), .A2(n1620), .Z(n1400) );
  and2 U1554 ( .A1(c), .A2(a), .Z(n1394) );
  and2 U1555 ( .A1(n1395), .A2(m), .Z(n1397) );
  and2 U1556 ( .A1(l), .A2(n1493), .Z(n1396) );
  or2 U1557 ( .A1(n1397), .A2(n1396), .Z(n1727) );
  inv1 U1558 ( .I(n1727), .ZN(n1398) );
  and2 U1559 ( .A1(n1156), .A2(n1398), .Z(n1399) );
  or2 U1560 ( .A1(n1400), .A2(n1399), .Z(n1401) );
  and2 U1564 ( .A1(n1628), .A2(n1254), .Z(n1407) );
  and2 U1565 ( .A1(n1630), .A2(n1673), .Z(n1406) );
  or2 U1566 ( .A1(n1406), .A2(n1407), .Z(n1408) );
  or2 U1568 ( .A1(n1161), .A2(n1409), .Z(n1800) );
  or2 U1570 ( .A1(n1522), .A2(l0), .Z(n1412) );
  inv1 U1571 ( .I(n1522), .ZN(n1410) );
  or2 U1572 ( .A1(n1410), .A2(h0), .Z(n1411) );
  and2 U1573 ( .A1(n1412), .A2(n1411), .Z(n1413) );
  and2 U1575 ( .A1(f0), .A2(n1607), .Z(n1414) );
  or2 U1576 ( .A1(n1415), .A2(n1414), .Z(n1419) );
  and2 U1577 ( .A1(n), .A2(n1601), .Z(n1417) );
  and2 U1578 ( .A1(g0), .A2(n1171), .Z(n1416) );
  or2 U1579 ( .A1(n1417), .A2(n1416), .Z(n1418) );
  or2 U1580 ( .A1(n1419), .A2(n1418), .Z(n1433) );
  or2 U1581 ( .A1(n1184), .A2(n1612), .Z(n1679) );
  inv1 U1582 ( .I(n1433), .ZN(n1672) );
  or2 U1583 ( .A1(n1672), .A2(n715), .Z(n1420) );
  or2 U1585 ( .A1(n1186), .A2(k), .Z(n1423) );
  or2 U1586 ( .A1(n1263), .A2(n1421), .Z(n1422) );
  and2 U1587 ( .A1(n1423), .A2(n1422), .Z(n1425) );
  and2 U1588 ( .A1(l), .A2(n1619), .Z(n1424) );
  or2 U1589 ( .A1(n1425), .A2(n1424), .Z(n1430) );
  and2 U1590 ( .A1(i), .A2(n1620), .Z(n1428) );
  and2 U1591 ( .A1(n1426), .A2(n1156), .Z(n1427) );
  or2 U1592 ( .A1(n1428), .A2(n1427), .Z(n1429) );
  or2 U1593 ( .A1(n1430), .A2(n1429), .Z(n1431) );
  and2 U1594 ( .A1(n1628), .A2(n1184), .Z(n1435) );
  and2 U1595 ( .A1(n1672), .A2(n1630), .Z(n1434) );
  inv1 U1601 ( .I(n1438), .ZN(n1490) );
  and2 U1602 ( .A1(m0), .A2(n1490), .Z(n1439) );
  and2 U1603 ( .A1(n1498), .A2(n1439), .Z(n1443) );
  inv1 U1604 ( .I(n1440), .ZN(n1496) );
  and2 U1605 ( .A1(l), .A2(n1496), .Z(n1441) );
  and2 U1606 ( .A1(n1498), .A2(n1441), .Z(n1442) );
  or2 U1607 ( .A1(n1443), .A2(n1442), .Z(n1448) );
  or2 U1608 ( .A1(n1186), .A2(n), .Z(n1446) );
  or2 U1609 ( .A1(n1156), .A2(n1444), .Z(n1445) );
  and2 U1610 ( .A1(n1263), .A2(n1446), .Z(n1447) );
  inv1 U1612 ( .I(n1450), .ZN(n1477) );
  and2 U1613 ( .A1(j0), .A2(n1477), .Z(n1452) );
  inv1 U1614 ( .I(n1188), .ZN(n1451) );
  and2 U1615 ( .A1(n1452), .A2(n1451), .Z(n1461) );
  and2 U1616 ( .A1(d), .A2(e), .Z(n1453) );
  or2 U1617 ( .A1(n1204), .A2(n1453), .Z(n1454) );
  inv1 U1618 ( .I(n1454), .ZN(n1457) );
  and2 U1619 ( .A1(o0), .A2(d), .Z(n1455) );
  and2 U1620 ( .A1(n1457), .A2(n1455), .Z(n1459) );
  and2 U1621 ( .A1(n1457), .A2(n1158), .Z(n1458) );
  or2 U1622 ( .A1(n1459), .A2(n1458), .Z(n1460) );
  and2 U1624 ( .A1(n1132), .A2(k0), .Z(n1462) );
  or2 U1626 ( .A1(n1480), .A2(n1463), .Z(n1464) );
  or2 U1630 ( .A1(n1467), .A2(n1466), .Z(n1468) );
  and2 U1631 ( .A1(n1658), .A2(n1468), .Z(n1472) );
  and2 U1634 ( .A1(n1469), .A2(n1470), .Z(n1471) );
  inv1 U1636 ( .I(n1178), .ZN(n1479) );
  and2 U1637 ( .A1(h0), .A2(n1159), .Z(n1473) );
  and2 U1638 ( .A1(n1479), .A2(n1473), .Z(n1476) );
  and2 U1639 ( .A1(n0), .A2(d), .Z(n1474) );
  and2 U1640 ( .A1(n1479), .A2(n1474), .Z(n1475) );
  or2 U1641 ( .A1(n1476), .A2(n1475), .Z(n1487) );
  and2 U1642 ( .A1(i0), .A2(n1477), .Z(n1478) );
  and2 U1643 ( .A1(n1479), .A2(n1478), .Z(n1481) );
  and2 U1645 ( .A1(j0), .A2(n1132), .Z(n1483) );
  and2 U1646 ( .A1(n1281), .A2(n1483), .Z(n1484) );
  or2 U1649 ( .A1(n1266), .A2(n1612), .Z(n1489) );
  or2 U1651 ( .A1(n1670), .A2(n715), .Z(n1488) );
  and2 U1652 ( .A1(n), .A2(n1490), .Z(n1491) );
  and2 U1653 ( .A1(n1498), .A2(n1491), .Z(n1501) );
  or2 U1654 ( .A1(n1186), .A2(m), .Z(n1492) );
  or2 U1655 ( .A1(n1156), .A2(n1492), .Z(n1495) );
  or2 U1656 ( .A1(n1263), .A2(n1493), .Z(n1494) );
  and2 U1657 ( .A1(n1495), .A2(n1494), .Z(n1500) );
  and2 U1658 ( .A1(k), .A2(n1496), .Z(n1497) );
  and2 U1659 ( .A1(n1498), .A2(n1497), .Z(n1499) );
  or2 U1660 ( .A1(n1500), .A2(n1197), .Z(n1504) );
  inv1 U1661 ( .I(n1504), .ZN(n1651) );
  or2 U1662 ( .A1(n1266), .A2(y), .Z(n1503) );
  or2 U1663 ( .A1(n1670), .A2(z), .Z(n1502) );
  inv1 U1666 ( .I(n1643), .ZN(n1506) );
  or2 U1667 ( .A1(n1506), .A2(n1218), .Z(n1653) );
  or2 U1669 ( .A1(n1508), .A2(n1507), .Z(n1669) );
  inv1 U1670 ( .I(n1669), .ZN(n1637) );
  or2 U1671 ( .A1(n1186), .A2(g), .Z(n1512) );
  or2 U1672 ( .A1(a), .A2(n1695), .Z(n1510) );
  or2 U1674 ( .A1(n1616), .A2(n1156), .Z(n1548) );
  or2 U1675 ( .A1(n1548), .A2(n2051), .Z(n1511) );
  and2 U1676 ( .A1(n1512), .A2(n1511), .Z(n1514) );
  and2 U1677 ( .A1(h), .A2(n1619), .Z(n1513) );
  or2 U1678 ( .A1(n1514), .A2(n1513), .Z(n1519) );
  and2 U1679 ( .A1(u), .A2(n1620), .Z(n1517) );
  and2 U1680 ( .A1(n1515), .A2(n1156), .Z(n1516) );
  or2 U1681 ( .A1(n1517), .A2(n1516), .Z(n1518) );
  or2 U1682 ( .A1(n1519), .A2(n1518), .Z(n1520) );
  inv1 U1683 ( .I(n1520), .ZN(n1910) );
  and2 U1684 ( .A1(b0), .A2(n1607), .Z(n1526) );
  inv1 U1685 ( .I(e), .ZN(n1521) );
  or2 U1686 ( .A1(a), .A2(n1521), .Z(n1523) );
  and2 U1689 ( .A1(d0), .A2(n1604), .Z(n1525) );
  or2 U1690 ( .A1(n1526), .A2(n1525), .Z(n1536) );
  and2 U1691 ( .A1(j), .A2(n1601), .Z(n1534) );
  and2 U1692 ( .A1(c0), .A2(n1171), .Z(n1532) );
  or2 U1694 ( .A1(a), .A2(n1528), .Z(n1529) );
  or2 U1695 ( .A1(n1530), .A2(n1529), .Z(n1531) );
  inv1 U1696 ( .I(n1531), .ZN(n1609) );
  or2 U1697 ( .A1(n1532), .A2(n1609), .Z(n1533) );
  or2 U1698 ( .A1(n1534), .A2(n1533), .Z(n1535) );
  or2 U1699 ( .A1(n1536), .A2(n1535), .Z(n1540) );
  and2 U1700 ( .A1(n1628), .A2(n1540), .Z(n1538) );
  inv1 U1701 ( .I(n1540), .ZN(n1541) );
  and2 U1702 ( .A1(n1630), .A2(n1541), .Z(n1537) );
  or2 U1703 ( .A1(n1538), .A2(n1537), .Z(n1539) );
  and2 U1704 ( .A1(n1910), .A2(n1539), .Z(n1546) );
  or2 U1705 ( .A1(n1540), .A2(n1612), .Z(n1543) );
  or2 U1706 ( .A1(n1541), .A2(n715), .Z(n1542) );
  and2 U1707 ( .A1(n1543), .A2(n1542), .Z(n1544) );
  or2 U1711 ( .A1(n1186), .A2(j), .Z(n1550) );
  or2 U1712 ( .A1(n1548), .A2(n1547), .Z(n1549) );
  and2 U1713 ( .A1(n1550), .A2(n1549), .Z(n1554) );
  and2 U1714 ( .A1(k), .A2(n1619), .Z(n1552) );
  and2 U1715 ( .A1(h), .A2(n1620), .Z(n1551) );
  or2 U1716 ( .A1(n1552), .A2(n1551), .Z(n1553) );
  and2 U1720 ( .A1(n1281), .A2(n1213), .Z(n1556) );
  and2 U1722 ( .A1(m), .A2(n1601), .Z(n1560) );
  or2 U1724 ( .A1(n1558), .A2(n1609), .Z(n1559) );
  or2 U1725 ( .A1(n1560), .A2(n1559), .Z(n1561) );
  and2 U1727 ( .A1(n1628), .A2(n1208), .Z(n1564) );
  inv1 U1728 ( .I(n1566), .ZN(n1567) );
  and2 U1729 ( .A1(n1630), .A2(n1567), .Z(n1563) );
  or2 U1730 ( .A1(n1564), .A2(n1563), .Z(n1565) );
  and2 U1731 ( .A1(n1710), .A2(n1565), .Z(n1571) );
  or2 U1732 ( .A1(n1208), .A2(n1612), .Z(n1569) );
  or2 U1733 ( .A1(n1567), .A2(n715), .Z(n1568) );
  and2 U1734 ( .A1(n1569), .A2(n1568), .Z(n1570) );
  inv1 U1736 ( .I(n1880), .ZN(n1638) );
  or2 U1738 ( .A1(n1186), .A2(h), .Z(n1573) );
  or2 U1739 ( .A1(n1249), .A2(n2050), .Z(n1572) );
  and2 U1740 ( .A1(n1573), .A2(n1572), .Z(n1575) );
  and2 U1741 ( .A1(i), .A2(n1619), .Z(n1574) );
  or2 U1742 ( .A1(n1575), .A2(n1574), .Z(n1582) );
  and2 U1743 ( .A1(v), .A2(n1620), .Z(n1580) );
  and2 U1744 ( .A1(h), .A2(i), .Z(n1577) );
  or2 U1745 ( .A1(n1577), .A2(n1576), .Z(n1578) );
  and2 U1746 ( .A1(n1156), .A2(n1578), .Z(n1579) );
  or2 U1747 ( .A1(n1580), .A2(n1579), .Z(n1581) );
  or2 U1748 ( .A1(n1582), .A2(n1581), .Z(n1583) );
  inv1 U1749 ( .I(n1583), .ZN(n1731) );
  and2 U1750 ( .A1(c0), .A2(n1607), .Z(n1585) );
  and2 U1751 ( .A1(e0), .A2(n1604), .Z(n1584) );
  or2 U1752 ( .A1(n1585), .A2(n1584), .Z(n1590) );
  and2 U1753 ( .A1(k), .A2(n1601), .Z(n1588) );
  and2 U1754 ( .A1(d0), .A2(n1171), .Z(n1586) );
  or2 U1755 ( .A1(n1586), .A2(n1609), .Z(n1587) );
  or2 U1756 ( .A1(n1588), .A2(n1587), .Z(n1589) );
  or2 U1757 ( .A1(n1590), .A2(n1589), .Z(n1594) );
  and2 U1758 ( .A1(n1628), .A2(n1594), .Z(n1592) );
  inv1 U1759 ( .I(n1594), .ZN(n1595) );
  and2 U1760 ( .A1(n1630), .A2(n1595), .Z(n1591) );
  or2 U1761 ( .A1(n1592), .A2(n1591), .Z(n1593) );
  and2 U1762 ( .A1(n1731), .A2(n1593), .Z(n1600) );
  or2 U1763 ( .A1(n1594), .A2(n1612), .Z(n1597) );
  or2 U1764 ( .A1(n1595), .A2(n715), .Z(n1596) );
  and2 U1765 ( .A1(n1597), .A2(n1596), .Z(n1598) );
  or2 U1768 ( .A1(n1600), .A2(n1757), .Z(n1733) );
  and2 U1769 ( .A1(e0), .A2(n1171), .Z(n1603) );
  or2 U1771 ( .A1(n1603), .A2(n1602), .Z(n1606) );
  or2 U1776 ( .A1(n1611), .A2(n1610), .Z(n1627) );
  or2 U1777 ( .A1(n1245), .A2(n1612), .Z(n1614) );
  inv1 U1778 ( .I(n1627), .ZN(n1629) );
  or2 U1779 ( .A1(n1629), .A2(n715), .Z(n1613) );
  and2 U1780 ( .A1(n1614), .A2(n1613), .Z(n1626) );
  or2 U1781 ( .A1(n1186), .A2(i), .Z(n1615) );
  or2 U1782 ( .A1(n1615), .A2(n1156), .Z(n1618) );
  or2 U1783 ( .A1(n1249), .A2(n2049), .Z(n1617) );
  and2 U1784 ( .A1(n1618), .A2(n1617), .Z(n1624) );
  and2 U1785 ( .A1(j), .A2(n1619), .Z(n1622) );
  and2 U1786 ( .A1(g), .A2(n1620), .Z(n1621) );
  or2 U1787 ( .A1(n1622), .A2(n1621), .Z(n1623) );
  or2 U1788 ( .A1(n1624), .A2(n1623), .Z(n1625) );
  and2 U1789 ( .A1(n1628), .A2(n1245), .Z(n1632) );
  and2 U1790 ( .A1(n1630), .A2(n1629), .Z(n1631) );
  or2 U1791 ( .A1(n1632), .A2(n1631), .Z(n1633) );
  and2 U1792 ( .A1(n1248), .A2(n1633), .Z(n1634) );
  or2 U1793 ( .A1(n1212), .A2(n1634), .Z(n1740) );
  and2 U1797 ( .A1(n1637), .A2(n1886), .Z(d1) );
  inv1 U1798 ( .I(n1913), .ZN(n1915) );
  inv1 U1799 ( .I(n1733), .ZN(n1735) );
  inv1 U1800 ( .I(n1740), .ZN(n1742) );
  and2 U1801 ( .A1(n1742), .A2(n1638), .Z(n1639) );
  and2 U1802 ( .A1(n1915), .A2(n1640), .Z(n1642) );
  or2 U1803 ( .A1(n1642), .A2(n1641), .Z(n1755) );
  inv1 U1804 ( .I(n1262), .ZN(n1802) );
  and2 U1811 ( .A1(n1886), .A2(n1754), .Z(n1648) );
  or2 U1812 ( .A1(n1198), .A2(n1648), .Z(e1) );
  or2 U1813 ( .A1(a), .A2(c), .Z(n1650) );
  inv1 U1814 ( .I(a0), .ZN(n1976) );
  or2 U1815 ( .A1(n1205), .A2(n1976), .Z(n1649) );
  or2 U1816 ( .A1(n1650), .A2(n1649), .Z(n1911) );
  inv1 U1817 ( .I(v0), .ZN(n1962) );
  or2 U1818 ( .A1(n1911), .A2(n1962), .Z(n1798) );
  and2 U1819 ( .A1(n1153), .A2(n1798), .Z(n1668) );
  or2 U1820 ( .A1(n1798), .A2(n1651), .Z(n1654) );
  inv1 U1821 ( .I(n1654), .ZN(n1652) );
  and2 U1822 ( .A1(n1246), .A2(n1652), .Z(n1657) );
  inv1 U1823 ( .I(n1246), .ZN(n1655) );
  and2 U1824 ( .A1(n1655), .A2(n1654), .Z(n1656) );
  or2 U1825 ( .A1(n1657), .A2(n1656), .Z(n1834) );
  or2 U1827 ( .A1(n1798), .A2(n1658), .Z(n1661) );
  inv1 U1828 ( .I(n1661), .ZN(n1659) );
  inv1 U1830 ( .I(n1660), .ZN(n1662) );
  and2 U1831 ( .A1(n1662), .A2(n1661), .Z(n1663) );
  inv1 U1838 ( .I(n1798), .ZN(n1881) );
  or2 U1839 ( .A1(n1670), .A2(n1671), .Z(n1676) );
  or2 U1840 ( .A1(n1672), .A2(x), .Z(n1674) );
  or2 U1841 ( .A1(n1674), .A2(n1231), .Z(n1675) );
  or2 U1842 ( .A1(n1676), .A2(n1675), .Z(n1684) );
  or2 U1843 ( .A1(n1254), .A2(n1679), .Z(n1681) );
  or2 U1844 ( .A1(n1682), .A2(n1681), .Z(n1683) );
  and2 U1845 ( .A1(n1684), .A2(n1683), .Z(n1685) );
  or2 U1846 ( .A1(n1685), .A2(n1798), .Z(n1867) );
  or2 U1849 ( .A1(n1829), .A2(a), .Z(n1692) );
  inv1 U1850 ( .I(n1688), .ZN(n1689) );
  and2 U1851 ( .A1(n1905), .A2(n1689), .Z(n1690) );
  or2 U1852 ( .A1(n1690), .A2(n2059), .Z(n1691) );
  and2 U1853 ( .A1(n1692), .A2(n1691), .Z(n1693) );
  or2 U1854 ( .A1(n1693), .A2(n741), .Z(g1) );
  and2 U1855 ( .A1(f), .A2(b), .Z(n1694) );
  and2 U1856 ( .A1(n1695), .A2(n1694), .Z(n1697) );
  or2 U1857 ( .A1(n1697), .A2(n2059), .Z(n1965) );
  or2 U1858 ( .A1(n1965), .A2(n2046), .Z(n1941) );
  inv1 U1859 ( .I(n1703), .ZN(n1698) );
  and2 U1860 ( .A1(u0), .A2(n1698), .Z(n1700) );
  inv1 U1861 ( .I(u0), .ZN(n1868) );
  and2 U1862 ( .A1(n1868), .A2(n1703), .Z(n1699) );
  or2 U1863 ( .A1(n1700), .A2(n1699), .Z(n1701) );
  and2 U1864 ( .A1(n1941), .A2(n1701), .Z(n1709) );
  inv1 U1865 ( .I(n1941), .ZN(n1856) );
  and2 U1866 ( .A1(n665), .A2(n1856), .Z(n1707) );
  inv1 U1867 ( .I(n1702), .ZN(n1853) );
  or2 U1868 ( .A1(n1703), .A2(n1853), .Z(n1705) );
  or2 U1869 ( .A1(n1937), .A2(n667), .Z(n1704) );
  and2 U1870 ( .A1(n1705), .A2(n1704), .Z(n1706) );
  and2 U1871 ( .A1(n1707), .A2(n1706), .Z(n1708) );
  or2 U1872 ( .A1(n1709), .A2(n1708), .Z(h1) );
  or2 U1873 ( .A1(n1710), .A2(n1798), .Z(n1713) );
  inv1 U1874 ( .I(n1713), .ZN(n1711) );
  and2 U1876 ( .A1(n1225), .A2(n1713), .Z(n1714) );
  and2 U1879 ( .A1(n1829), .A2(n1878), .Z(n1717) );
  or2 U1880 ( .A1(n1141), .A2(n1716), .Z(n1718) );
  and2 U1882 ( .A1(n614), .A2(n1856), .Z(n1723) );
  or2 U1883 ( .A1(n1719), .A2(n136), .Z(n1721) );
  or2 U1884 ( .A1(n1937), .A2(n616), .Z(n1720) );
  and2 U1885 ( .A1(n1721), .A2(n1720), .Z(n1722) );
  inv1 U1887 ( .I(n1775), .ZN(n1726) );
  and2 U1888 ( .A1(n550), .A2(n1726), .Z(n1786) );
  and2 U1889 ( .A1(n), .A2(n1727), .Z(n1729) );
  or2 U1890 ( .A1(n1729), .A2(n1728), .Z(n1784) );
  or2 U1891 ( .A1(n1869), .A2(n1730), .Z(n1749) );
  inv1 U1892 ( .I(n1749), .ZN(n1747) );
  or2 U1893 ( .A1(n1911), .A2(n1731), .Z(n1734) );
  inv1 U1894 ( .I(n1734), .ZN(n1732) );
  and2 U1895 ( .A1(n1733), .A2(n1732), .Z(n1737) );
  and2 U1896 ( .A1(n1735), .A2(n1734), .Z(n1736) );
  or2 U1900 ( .A1(n1798), .A2(n1248), .Z(n1741) );
  inv1 U1901 ( .I(n1741), .ZN(n1739) );
  or2 U1906 ( .A1(n1875), .A2(n1878), .Z(n1745) );
  or2 U1908 ( .A1(n1747), .A2(n1748), .Z(n1751) );
  inv1 U1909 ( .I(n1748), .ZN(n1907) );
  or2 U1910 ( .A1(n1749), .A2(n1907), .Z(n1750) );
  and2 U1911 ( .A1(n1751), .A2(n1750), .Z(n1752) );
  or2 U1912 ( .A1(n1752), .A2(n1868), .Z(n1778) );
  inv1 U1913 ( .I(n1778), .ZN(n1773) );
  and2 U1914 ( .A1(n1886), .A2(n1798), .Z(n1753) );
  and2 U1915 ( .A1(n1754), .A2(n1753), .Z(n1756) );
  or2 U1916 ( .A1(n1755), .A2(n1756), .Z(n1889) );
  and2 U1917 ( .A1(n1757), .A2(n1911), .Z(n1768) );
  and2 U1918 ( .A1(n1199), .A2(n1880), .Z(n1763) );
  and2 U1919 ( .A1(n1758), .A2(n1180), .Z(n1761) );
  and2 U1920 ( .A1(n1180), .A2(n1280), .Z(n1759) );
  or2 U1921 ( .A1(n1759), .A2(n1140), .Z(n1760) );
  or2 U1928 ( .A1(n1768), .A2(n1864), .Z(n1908) );
  inv1 U1929 ( .I(n1908), .ZN(n1769) );
  and2 U1930 ( .A1(n1889), .A2(n1769), .Z(n1772) );
  inv1 U1931 ( .I(n1889), .ZN(n1770) );
  and2 U1932 ( .A1(n1770), .A2(n1908), .Z(n1771) );
  or2 U1933 ( .A1(n1772), .A2(n1771), .Z(n1776) );
  or2 U1934 ( .A1(n1773), .A2(n1776), .Z(n1774) );
  and2 U1935 ( .A1(n1775), .A2(n1774), .Z(n1780) );
  inv1 U1936 ( .I(n1776), .ZN(n1777) );
  or2 U1937 ( .A1(n1778), .A2(n1777), .Z(n1779) );
  and2 U1938 ( .A1(n1780), .A2(n1779), .Z(n1782) );
  or2 U1939 ( .A1(n1782), .A2(n1781), .Z(n1783) );
  and2 U1940 ( .A1(n1784), .A2(n1783), .Z(n1785) );
  or2 U1941 ( .A1(n1786), .A2(n1785), .Z(j1) );
  or2 U1942 ( .A1(n1798), .A2(n1194), .Z(n1789) );
  inv1 U1943 ( .I(n1789), .ZN(n1787) );
  and2 U1944 ( .A1(n1280), .A2(n1787), .Z(n1791) );
  and2 U1945 ( .A1(n1230), .A2(n1789), .Z(n1790) );
  or2 U1946 ( .A1(n1791), .A2(n1790), .Z(n1809) );
  or2 U1947 ( .A1(n1809), .A2(n1853), .Z(n1792) );
  and2 U1948 ( .A1(n1856), .A2(n1792), .Z(n1796) );
  or2 U1949 ( .A1(n1937), .A2(n461), .Z(n1794) );
  or2 U1950 ( .A1(n377), .A2(n493), .Z(n1793) );
  and2 U1951 ( .A1(n1794), .A2(n1793), .Z(n1795) );
  and2 U1952 ( .A1(n1796), .A2(n1795), .Z(n1828) );
  and2 U1953 ( .A1(n1161), .A2(n1798), .Z(n1806) );
  or2 U1954 ( .A1(n1798), .A2(n1797), .Z(n1801) );
  inv1 U1955 ( .I(n1801), .ZN(n1799) );
  and2 U1956 ( .A1(n1800), .A2(n1799), .Z(n1804) );
  and2 U1957 ( .A1(n1802), .A2(n1801), .Z(n1803) );
  or2 U1958 ( .A1(n1804), .A2(n1803), .Z(n1854) );
  inv1 U1961 ( .I(n1809), .ZN(n1807) );
  and2 U1962 ( .A1(n1808), .A2(n1807), .Z(n1812) );
  inv1 U1963 ( .I(n1808), .ZN(n1810) );
  and2 U1964 ( .A1(n1810), .A2(n1809), .Z(n1811) );
  or2 U1965 ( .A1(n1812), .A2(n1811), .Z(n1826) );
  inv1 U1966 ( .I(n1834), .ZN(n1813) );
  and2 U1967 ( .A1(n1813), .A2(n1814), .Z(n1817) );
  inv1 U1968 ( .I(n1814), .ZN(n1815) );
  and2 U1969 ( .A1(n1834), .A2(n1815), .Z(n1816) );
  or2 U1970 ( .A1(n1817), .A2(n1816), .Z(n1831) );
  inv1 U1972 ( .I(n1854), .ZN(n1818) );
  and2 U1973 ( .A1(f1), .A2(n1818), .Z(n1821) );
  inv1 U1974 ( .I(f1), .ZN(n1819) );
  and2 U1977 ( .A1(n1822), .A2(n1846), .Z(n1824) );
  or2 U1980 ( .A1(n1824), .A2(n1847), .Z(n1825) );
  or2 U1983 ( .A1(n1829), .A2(n1905), .Z(n1842) );
  inv1 U1984 ( .I(n1842), .ZN(n1830) );
  inv1 U1986 ( .I(n1831), .ZN(n1845) );
  or2 U1987 ( .A1(n1845), .A2(n1847), .Z(n1832) );
  or2 U1989 ( .A1(n1834), .A2(n1853), .Z(n1835) );
  and2 U1990 ( .A1(n1856), .A2(n1835), .Z(n1839) );
  or2 U1991 ( .A1(n1937), .A2(n401), .Z(n1837) );
  or2 U1992 ( .A1(n377), .A2(n435), .Z(n1836) );
  and2 U1993 ( .A1(n1837), .A2(n1836), .Z(n1838) );
  and2 U1994 ( .A1(n1839), .A2(n1838), .Z(n1840) );
  or2 U1995 ( .A1(n1841), .A2(n1840), .Z(l1) );
  or2 U1996 ( .A1(n1842), .A2(n1845), .Z(n1843) );
  inv1 U1997 ( .I(n1843), .ZN(n1844) );
  or2 U1998 ( .A1(n1844), .A2(n1846), .Z(n1852) );
  and2 U1999 ( .A1(n2046), .A2(n1845), .Z(n1850) );
  inv1 U2000 ( .I(n1846), .ZN(n1848) );
  or2 U2001 ( .A1(n1848), .A2(n1847), .Z(n1849) );
  or2 U2002 ( .A1(n1850), .A2(n1849), .Z(n1851) );
  or2 U2004 ( .A1(n1854), .A2(n1853), .Z(n1855) );
  and2 U2005 ( .A1(n1856), .A2(n1855), .Z(n1860) );
  or2 U2006 ( .A1(n1937), .A2(n342), .Z(n1858) );
  or2 U2007 ( .A1(n377), .A2(n376), .Z(n1857) );
  and2 U2008 ( .A1(n1858), .A2(n1857), .Z(n1859) );
  and2 U2009 ( .A1(n1860), .A2(n1859), .Z(n1861) );
  and2 U2013 ( .A1(n1866), .A2(n1867), .Z(n1869) );
  or2 U2014 ( .A1(n1150), .A2(n1154), .Z(n1874) );
  inv1 U2015 ( .I(n1264), .ZN(n1877) );
  inv1 U2017 ( .I(n1903), .ZN(n1872) );
  or2 U2018 ( .A1(n1873), .A2(n1872), .Z(n1895) );
  inv1 U2019 ( .I(n1895), .ZN(n1964) );
  and2 U2020 ( .A1(n1874), .A2(n1875), .Z(n1876) );
  and2 U2022 ( .A1(n1243), .A2(n1180), .Z(n1879) );
  inv1 U2026 ( .I(n1946), .ZN(n1978) );
  and2 U2027 ( .A1(u0), .A2(n1886), .Z(n1887) );
  and2 U2028 ( .A1(n1888), .A2(n1887), .Z(n1890) );
  inv1 U2031 ( .I(n1891), .ZN(n1892) );
  inv1 U2034 ( .I(n132), .ZN(n1924) );
  and2 U2035 ( .A1(n2050), .A2(n1924), .Z(n1897) );
  and2 U2036 ( .A1(n275), .A2(n1925), .Z(n1896) );
  or2 U2037 ( .A1(n1897), .A2(n1896), .Z(n1901) );
  and2 U2038 ( .A1(n152), .A2(n1898), .Z(n1899) );
  or2 U2039 ( .A1(n1899), .A2(n1941), .Z(n1900) );
  or2 U2040 ( .A1(n1901), .A2(n1900), .Z(n1969) );
  inv1 U2041 ( .I(n1948), .ZN(n1945) );
  or2 U2042 ( .A1(n1903), .A2(n1978), .Z(n1904) );
  and2 U2045 ( .A1(u0), .A2(n1907), .Z(n1909) );
  or2 U2046 ( .A1(n1911), .A2(n1910), .Z(n1914) );
  inv1 U2047 ( .I(n1914), .ZN(n1912) );
  and2 U2048 ( .A1(n1913), .A2(n1912), .Z(n1917) );
  and2 U2049 ( .A1(n1915), .A2(n1914), .Z(n1916) );
  or2 U2050 ( .A1(n1917), .A2(n1916), .Z(n1919) );
  inv1 U2051 ( .I(n1919), .ZN(n1928) );
  and2 U2052 ( .A1(n1918), .A2(n1928), .Z(n1922) );
  inv1 U2053 ( .I(n1918), .ZN(n1920) );
  and2 U2059 ( .A1(n2051), .A2(n1924), .Z(n1927) );
  and2 U2060 ( .A1(n157), .A2(n1925), .Z(n1926) );
  or2 U2061 ( .A1(n1927), .A2(n1926), .Z(n1931) );
  and2 U2062 ( .A1(n152), .A2(n1928), .Z(n1929) );
  or2 U2063 ( .A1(n1929), .A2(n1941), .Z(n1930) );
  or2 U2064 ( .A1(n1931), .A2(n1930), .Z(n1960) );
  inv1 U2065 ( .I(n1960), .ZN(n1934) );
  or2 U2068 ( .A1(n1936), .A2(n1935), .Z(n2052) );
  or2 U2069 ( .A1(i), .A2(n132), .Z(n1939) );
  or2 U2070 ( .A1(n86), .A2(n1937), .Z(n1938) );
  and2 U2071 ( .A1(n1939), .A2(n1938), .Z(n1944) );
  or2 U2072 ( .A1(n1940), .A2(n136), .Z(n1942) );
  and2 U2073 ( .A1(n1942), .A2(n1856), .Z(n1943) );
  and2 U2074 ( .A1(n1944), .A2(n1943), .Z(n1979) );
  and2 U2075 ( .A1(n1945), .A2(n2046), .Z(n1947) );
  or2 U2076 ( .A1(n1265), .A2(n1947), .Z(n1977) );
  or2 U2079 ( .A1(n1278), .A2(n1980), .Z(n1950) );
  and2 U2080 ( .A1(n1977), .A2(n1950), .Z(n1951) );
  or2 U2081 ( .A1(n1979), .A2(n1951), .Z(p1) );
  or2 U2082 ( .A1(h1), .A2(i1), .Z(n1953) );
  or2 U2083 ( .A1(k1), .A2(l1), .Z(n1952) );
  or2 U2084 ( .A1(n1953), .A2(n1952), .Z(n1957) );
  or2 U2085 ( .A1(m1), .A2(p1), .Z(n1955) );
  or2 U2086 ( .A1(o1), .A2(n1), .Z(n1954) );
  or2 U2087 ( .A1(n1955), .A2(n1954), .Z(n1956) );
  or2 U2088 ( .A1(n1957), .A2(n1956), .Z(q1) );
  inv1 U2089 ( .I(q1), .ZN(n1958) );
  or2 U2090 ( .A1(n1958), .A2(n1976), .Z(n1975) );
  and2 U2091 ( .A1(n1960), .A2(n1959), .Z(n1961) );
  and2 U2092 ( .A1(n1962), .A2(n1961), .Z(n1973) );
  and2 U2093 ( .A1(n1964), .A2(n1963), .Z(n1967) );
  inv1 U2094 ( .I(n1965), .ZN(n1966) );
  or2 U2095 ( .A1(n1967), .A2(n1966), .Z(n1968) );
  and2 U2096 ( .A1(n1969), .A2(n1968), .Z(n1970) );
  and2 U2097 ( .A1(n1971), .A2(n1970), .Z(n1972) );
  and2 U2098 ( .A1(n1973), .A2(n1972), .Z(n1974) );
  or2 U2099 ( .A1(n1975), .A2(n1974), .Z(r1) );
  or2 U2100 ( .A1(n1976), .A2(v0), .Z(n1994) );
  inv1 U2101 ( .I(n1994), .ZN(n1993) );
  or2 U2103 ( .A1(n1978), .A2(n1979), .Z(n1981) );
  inv1 U2106 ( .I(i1), .ZN(n1982) );
  or2 U2107 ( .A1(n1983), .A2(n1982), .Z(n1984) );
  inv1 U2111 ( .I(x0), .ZN(n1989) );
  or2 U2115 ( .A1(n1241), .A2(n1162), .Z(n2032) );
  inv1 U2121 ( .I(n2032), .ZN(n2030) );
  inv1 U2124 ( .I(m1), .ZN(n2001) );
  inv1 U2126 ( .I(h1), .ZN(n2002) );
  inv1 U2129 ( .I(l1), .ZN(n2005) );
  and2 U2130 ( .A1(n2005), .A2(k1), .Z(n2008) );
  and2 U2132 ( .A1(l1), .A2(n2006), .Z(n2007) );
  inv1 U2136 ( .I(n2010), .ZN(n2012) );
  inv1 U2141 ( .I(n2019), .ZN(n2020) );
  or2 U2142 ( .A1(n2020), .A2(n2027), .Z(n2021) );
  or2 U2147 ( .A1(n2031), .A2(n2030), .Z(n2035) );
  or2 U2149 ( .A1(n2033), .A2(n2032), .Z(n2034) );
  and2 U2150 ( .A1(n2035), .A2(n2034), .Z(t1) );
  and2f U1150 ( .A1(n1829), .A2(n1878), .Z(n1141) );
  or2f U1151 ( .A1(n1644), .A2(n1153), .Z(n1645) );
  inv1f U1152 ( .I(n1883), .ZN(n1234) );
  or2f U1153 ( .A1(n1646), .A2(n1161), .Z(n1647) );
  inv1f U1155 ( .I(n1405), .ZN(n1161) );
  inv1f U1156 ( .I(n1371), .ZN(n1171) );
  and2 U1157 ( .A1(f0), .A2(n1171), .Z(n1558) );
  inv1f U1161 ( .I(n1599), .ZN(n1757) );
  inv1f U1162 ( .I(n182), .ZN(n2042) );
  inv1f U1164 ( .I(n1509), .ZN(n1498) );
  and2f U1165 ( .A1(n1510), .A2(n1509), .Z(n1616) );
  or2f U1166 ( .A1(n1440), .A2(n1509), .Z(n1393) );
  inv1f U1171 ( .I(n1545), .ZN(n1641) );
  inv1 U1173 ( .I(n1393), .ZN(n1620) );
  and2 U1174 ( .A1(n1819), .A2(n1854), .Z(n1820) );
  and2 U1175 ( .A1(f0), .A2(n1604), .Z(n1605) );
  or2 U1176 ( .A1(d), .A2(n1370), .Z(n1450) );
  inv1 U1177 ( .I(n1555), .ZN(n1710) );
  and2 U1178 ( .A1(n1194), .A2(n1436), .Z(n1437) );
  or2 U1185 ( .A1(n1636), .A2(n1635), .Z(n1730) );
  and2 U1186 ( .A1(n1660), .A2(n1659), .Z(n1664) );
  or2 U1190 ( .A1(n1905), .A2(n1892), .Z(n1168) );
  inv1 U1191 ( .I(n1984), .ZN(n1241) );
  or2 U1198 ( .A1(n1544), .A2(n1910), .Z(n1545) );
  and2 U1199 ( .A1(n1723), .A2(n1722), .Z(n1724) );
  and2 U1202 ( .A1(n2046), .A2(n1831), .Z(n1822) );
  or2f U1204 ( .A1(n1527), .A2(a), .Z(n1365) );
  inv1 U1205 ( .I(n2041), .ZN(n2057) );
  inv1 U1206 ( .I(n2057), .ZN(n2058) );
  or2f U1207 ( .A1(n1165), .A2(n2059), .Z(n1509) );
  and2f U1208 ( .A1(n1524), .A2(n1281), .Z(n1604) );
  and2f U1210 ( .A1(n1281), .A2(n1462), .Z(n1463) );
  and2f U1211 ( .A1(n1281), .A2(n1413), .Z(n1415) );
  inv1f U1214 ( .I(n1678), .ZN(n1671) );
  or2f U1217 ( .A1(n1205), .A2(n1160), .Z(n1188) );
  or2f U1218 ( .A1(n1205), .A2(n2059), .Z(n1204) );
  and2f U1219 ( .A1(n2046), .A2(n1948), .Z(n1949) );
  or2f U1220 ( .A1(n1755), .A2(n1135), .Z(n1948) );
  or2 U1221 ( .A1(n1830), .A2(n1831), .Z(n1833) );
  inv1 U1222 ( .I(n1157), .ZN(n1281) );
  and2 U1231 ( .A1(n1202), .A2(n1192), .Z(n1157) );
  inv1 U1236 ( .I(n1387), .ZN(n1263) );
  or2 U1239 ( .A1(n1379), .A2(n1378), .Z(n1254) );
  or2 U1241 ( .A1(n2042), .A2(n2041), .Z(n104) );
  or2 U1242 ( .A1(n1225), .A2(n1196), .Z(n1195) );
  inv1 U1243 ( .I(n1738), .ZN(n1898) );
  inv1 U1244 ( .I(k1), .ZN(n2006) );
  and2 U1247 ( .A1(n1628), .A2(n1678), .Z(n1467) );
  and2 U1253 ( .A1(n1369), .A2(n1202), .Z(n1601) );
  or2 U1256 ( .A1(n1505), .A2(n1504), .Z(n1643) );
  inv1 U1260 ( .I(n1268), .ZN(n1712) );
  and2 U1261 ( .A1(n1226), .A2(n1227), .Z(n1173) );
  inv1 U1262 ( .I(n1932), .ZN(n1963) );
  or2 U1265 ( .A1(n1806), .A2(n1805), .Z(n1808) );
  and2 U1266 ( .A1(n1149), .A2(n1969), .Z(n1148) );
  inv1 U1270 ( .I(n1902), .ZN(n1149) );
  inv1 U1274 ( .I(n2011), .ZN(n2009) );
  or2 U1275 ( .A1(n1282), .A2(n1437), .Z(n1788) );
  or2 U1276 ( .A1(n1217), .A2(n1282), .Z(n1754) );
  inv1 U1277 ( .I(n1730), .ZN(n1886) );
  and2 U1278 ( .A1(n1143), .A2(n1798), .Z(n1666) );
  or2 U1279 ( .A1(n1949), .A2(n1965), .Z(n1980) );
  or2 U1280 ( .A1(n2026), .A2(n1998), .Z(n1258) );
  or2 U1285 ( .A1(n1725), .A2(n1724), .Z(i1) );
  and2 U1286 ( .A1(n1941), .A2(n1718), .Z(n1725) );
  and2 U1293 ( .A1(n1833), .A2(n1832), .Z(n1841) );
  or2 U1294 ( .A1(n1935), .A2(n1936), .Z(o1) );
  inv1f U1295 ( .I(b), .ZN(n1205) );
  and2f U1297 ( .A1(n1527), .A2(n1521), .Z(n1530) );
  or2 U1298 ( .A1(a), .A2(n1527), .Z(n1522) );
  or2 U1299 ( .A1(n1372), .A2(n1527), .Z(n1482) );
  or2 U1300 ( .A1(n1133), .A2(n1527), .Z(n1132) );
  inv1f U1301 ( .I(f), .ZN(n1527) );
  and2f U1302 ( .A1(g0), .A2(n1607), .Z(n1368) );
  and2 U1305 ( .A1(e0), .A2(n1607), .Z(n1557) );
  and2 U1306 ( .A1(n1607), .A2(d0), .Z(n1608) );
  inv1f U1307 ( .I(n1364), .ZN(n1607) );
  inv1f U1309 ( .I(a), .ZN(n2059) );
  inv1 U1311 ( .I(a), .ZN(n2060) );
  or2f U1313 ( .A1(n1384), .A2(n1186), .Z(n1385) );
  and2f U1314 ( .A1(c), .A2(n1175), .Z(n1186) );
  inv1 U1315 ( .I(n1677), .ZN(n1670) );
  inv1 U1316 ( .I(n1719), .ZN(n1878) );
  or2 U1318 ( .A1(n1715), .A2(n1714), .Z(n1719) );
  or2 U1319 ( .A1(n1465), .A2(n1464), .Z(n1257) );
  or2 U1320 ( .A1(n1404), .A2(n1797), .Z(n1405) );
  inv1 U1321 ( .I(n1647), .ZN(n1758) );
  inv1 U1323 ( .I(n2056), .ZN(n1985) );
  or2f U1325 ( .A1(n1438), .A2(n1509), .Z(n1390) );
  or2 U1330 ( .A1(n1162), .A2(n1989), .Z(n1235) );
  and2f U1331 ( .A1(n1987), .A2(n1988), .Z(n1162) );
  or2f U1380 ( .A1(n1210), .A2(n1211), .Z(n1209) );
  and2f U1413 ( .A1(n1763), .A2(n1762), .Z(n1766) );
  or2f U1416 ( .A1(n1761), .A2(n1760), .Z(n1762) );
  or2f U1428 ( .A1(n1188), .A2(n1450), .Z(n1371) );
  inv1f U1510 ( .I(n2027), .ZN(n2015) );
  inv1f U1511 ( .I(n1449), .ZN(n1658) );
  and2f U1513 ( .A1(n1214), .A2(n1215), .Z(n2056) );
  and2f U1517 ( .A1(n1971), .A2(n1148), .Z(n1255) );
  or2f U1518 ( .A1(n1879), .A2(n1228), .Z(n1226) );
  and2f U1519 ( .A1(n1647), .A2(n1230), .Z(n1229) );
  inv1f U1522 ( .I(n1403), .ZN(n1797) );
  or2f U1523 ( .A1(n1402), .A2(n1401), .Z(n1403) );
  or2f U1526 ( .A1(n1386), .A2(n1385), .Z(n1387) );
  or2f U1529 ( .A1(n1768), .A2(n1222), .Z(n1918) );
  or2f U1530 ( .A1(n1909), .A2(n1864), .Z(n1222) );
  and2f U1535 ( .A1(n1269), .A2(n1880), .Z(n1268) );
  or2f U1540 ( .A1(n1557), .A2(n1556), .Z(n1562) );
  or2f U1541 ( .A1(n1999), .A2(n2030), .Z(n2000) );
  inv1f U1545 ( .I(n1940), .ZN(n1875) );
  and2f U1546 ( .A1(n1884), .A2(n1173), .Z(n1129) );
  and2f U1551 ( .A1(l), .A2(n1601), .Z(n1602) );
  and2f U1552 ( .A1(n1136), .A2(n1739), .Z(n1744) );
  or2f U1561 ( .A1(n1521), .A2(n1284), .Z(n1202) );
  and2f U1562 ( .A1(n1863), .A2(n1898), .Z(n1865) );
  or2f U1563 ( .A1(n1766), .A2(n1765), .Z(n1863) );
  and2f U1567 ( .A1(n1904), .A2(n1945), .Z(n1906) );
  or2f U1569 ( .A1(n1554), .A2(n1553), .Z(n1555) );
  or2f U1574 ( .A1(n1666), .A2(n1665), .Z(n1814) );
  or2f U1584 ( .A1(n2004), .A2(n2003), .Z(n2010) );
  and2f U1596 ( .A1(m1), .A2(n2002), .Z(n2003) );
  and2f U1597 ( .A1(u0), .A2(n1703), .Z(n1665) );
  inv1f U1598 ( .I(n1130), .ZN(n1) );
  and2f U1599 ( .A1(n1971), .A2(n1148), .Z(n1130) );
  and2f U1600 ( .A1(n1965), .A2(n1895), .Z(n1902) );
  and2f U1611 ( .A1(n1523), .A2(n1522), .Z(n1524) );
  and2f U1623 ( .A1(n1134), .A2(n1274), .Z(n1142) );
  and2f U1625 ( .A1(n1993), .A2(n1273), .Z(n1134) );
  or2f U1627 ( .A1(n1283), .A2(x0), .Z(n1274) );
  or2f U1628 ( .A1(n1733), .A2(n1136), .Z(n1635) );
  or2f U1629 ( .A1(n1546), .A2(n1641), .Z(n1913) );
  or2f U1632 ( .A1(n1756), .A2(n1890), .Z(n1135) );
  and2f U1633 ( .A1(n2010), .A2(n2009), .Z(n2014) );
  and2f U1635 ( .A1(n1826), .A2(n1825), .Z(n1827) );
  and2f U1644 ( .A1(f1), .A2(n1854), .Z(n1805) );
  and2f U1647 ( .A1(n2060), .A2(b), .Z(n1175) );
  inv1f U1648 ( .I(n1959), .ZN(n1936) );
  inv1f U1650 ( .I(n2031), .ZN(n2033) );
  or2f U1664 ( .A1(n1562), .A2(n1561), .Z(n1566) );
  and2f U1665 ( .A1(n1993), .A2(n1992), .Z(n1277) );
  and2f U1668 ( .A1(n1987), .A2(n1988), .Z(n1995) );
  or2f U1673 ( .A1(n1277), .A2(n1994), .Z(n2019) );
  or2f U1687 ( .A1(n1172), .A2(n1179), .Z(n1177) );
  inv1f U1688 ( .I(n1207), .ZN(n1179) );
  or2f U1693 ( .A1(n1609), .A2(n1608), .Z(n1610) );
  and2f U1708 ( .A1(n1991), .A2(n1142), .Z(n1276) );
  or2f U1709 ( .A1(n1800), .A2(n1788), .Z(n1508) );
  and2f U1710 ( .A1(u0), .A2(n1888), .Z(n1686) );
  inv1f U1717 ( .I(n1150), .ZN(n1888) );
  or2f U1718 ( .A1(n1435), .A2(n1434), .Z(n1436) );
  and2f U1719 ( .A1(n2015), .A2(n1139), .Z(n2029) );
  or2f U1721 ( .A1(n1922), .A2(n1921), .Z(n1932) );
  and2f U1723 ( .A1(n1920), .A2(n1919), .Z(n1921) );
  or2f U1726 ( .A1(n1746), .A2(n1745), .Z(n1748) );
  or2f U1735 ( .A1(n1898), .A2(n1869), .Z(n1746) );
  or2f U1737 ( .A1(n1598), .A2(n1731), .Z(n1599) );
  or2f U1766 ( .A1(n1737), .A2(n1736), .Z(n1738) );
  or2f U1767 ( .A1(n1997), .A2(n1996), .Z(n2025) );
  or2f U1770 ( .A1(n1486), .A2(n1487), .Z(n1677) );
  and2f U1772 ( .A1(n1802), .A2(n1645), .Z(n1646) );
  or2f U1773 ( .A1(n1485), .A2(n1484), .Z(n1486) );
  or2f U1774 ( .A1(n1481), .A2(n1480), .Z(n1485) );
  and2f U1775 ( .A1(n1503), .A2(n1502), .Z(n1505) );
  or2f U1794 ( .A1(n1894), .A2(n1893), .Z(n1971) );
  and2f U1795 ( .A1(n1964), .A2(n1891), .Z(n1894) );
  and2f U1796 ( .A1(n1167), .A2(n1168), .Z(n1893) );
  or2f U1805 ( .A1(n1235), .A2(n1241), .Z(n1991) );
  and2f U1806 ( .A1(n1993), .A2(n1992), .Z(n1999) );
  and2f U1807 ( .A1(n1712), .A2(n1711), .Z(n1715) );
  and2f U1808 ( .A1(n1988), .A2(n1986), .Z(n1983) );
  or2f U1809 ( .A1(n1981), .A2(n1980), .Z(n1988) );
  and2f U1810 ( .A1(n1884), .A2(n1173), .Z(n1885) );
  and2f U1826 ( .A1(n2001), .A2(h1), .Z(n2004) );
  or2f U1829 ( .A1(n1465), .A2(n1464), .Z(n1678) );
  or2f U1832 ( .A1(n1668), .A2(n1667), .Z(f1) );
  and2f U1833 ( .A1(n1834), .A2(n1814), .Z(n1667) );
  or2f U1834 ( .A1(n1862), .A2(n1861), .Z(m1) );
  and2f U1835 ( .A1(n1852), .A2(n1851), .Z(n1862) );
  or2f U1836 ( .A1(n1460), .A2(n1461), .Z(n1465) );
  or2f U1837 ( .A1(n1276), .A2(n2032), .Z(n1998) );
  or2f U1847 ( .A1(n1885), .A2(n1232), .Z(n1946) );
  and2f U1848 ( .A1(n1143), .A2(n1643), .Z(n1644) );
  or2f U1875 ( .A1(n1678), .A2(n1612), .Z(n1470) );
  inv1f U1877 ( .I(n1147), .ZN(s1) );
  or2f U1878 ( .A1(n1998), .A2(n1220), .Z(n2018) );
  or2f U1881 ( .A1(n1983), .A2(n1275), .Z(n1273) );
  or2f U1886 ( .A1(n1278), .A2(n1948), .Z(n1891) );
  or2f U1897 ( .A1(n1712), .A2(n1913), .Z(n1636) );
  or2f U1898 ( .A1(n2008), .A2(n2007), .Z(n2011) );
  or2f U1899 ( .A1(n1828), .A2(n1827), .Z(k1) );
  or2f U1902 ( .A1(n1821), .A2(n1820), .Z(n1846) );
  or2f U1903 ( .A1(n1151), .A2(n1472), .Z(n1660) );
  or2f U1904 ( .A1(n1664), .A2(n1663), .Z(n1703) );
  and2f U1905 ( .A1(n2027), .A2(n2026), .Z(n2028) );
  and2f U1907 ( .A1(n1871), .A2(n1877), .Z(n1873) );
  or2f U1922 ( .A1(n1864), .A2(n1170), .Z(n1871) );
  and2f U1923 ( .A1(n1797), .A2(n1408), .Z(n1409) );
  or2f U1924 ( .A1(n1996), .A2(n1997), .Z(n1139) );
  and2f U1925 ( .A1(o1), .A2(n1130), .Z(n1997) );
  or2f U1926 ( .A1(n1480), .A2(n1368), .Z(n1379) );
  and2f U1927 ( .A1(n2017), .A2(n1258), .Z(n1146) );
  or2f U1959 ( .A1(n1139), .A2(n2000), .Z(n2017) );
  and2f U1960 ( .A1(n1991), .A2(n1990), .Z(n1992) );
  and2f U1971 ( .A1(n1274), .A2(n1273), .Z(n1990) );
  and2f U1975 ( .A1(n1986), .A2(n1985), .Z(n1987) );
  or2f U1976 ( .A1(n1244), .A2(n1947), .Z(n1986) );
  and2f U1978 ( .A1(n1866), .A2(n1867), .Z(n1150) );
  or2f U1979 ( .A1(n1508), .A2(n1253), .Z(n1866) );
  or2f U1981 ( .A1(n1876), .A2(n1272), .Z(n1882) );
  inv1f U1982 ( .I(n1870), .ZN(n1272) );
  or2f U1985 ( .A1(n1432), .A2(n1194), .Z(n1180) );
  and2f U1988 ( .A1(n1679), .A2(n1420), .Z(n1432) );
  inv1f U2003 ( .I(n1139), .ZN(n2026) );
  or2f U2010 ( .A1(n1233), .A2(n1885), .Z(n1265) );
  and2f U2011 ( .A1(n1882), .A2(n1234), .Z(n1232) );
  and2f U2012 ( .A1(n1882), .A2(n1234), .Z(n1233) );
  inv1f U2016 ( .I(n1882), .ZN(n1884) );
  or2f U2021 ( .A1(n1653), .A2(n1660), .Z(n1507) );
  or2f U2023 ( .A1(n1671), .A2(n715), .Z(n1469) );
  or2f U2024 ( .A1(y), .A2(n1257), .Z(n1200) );
  inv1f U2025 ( .I(n1187), .ZN(n1996) );
  or2f U2029 ( .A1(n1255), .A2(n2052), .Z(n1187) );
  and2f U2030 ( .A1(n1261), .A2(n2017), .Z(n2016) );
  or2f U2032 ( .A1(n1923), .A2(n1963), .Z(n1959) );
  or2f U2033 ( .A1(n1906), .A2(n1905), .Z(n1923) );
  or2f U2043 ( .A1(n1864), .A2(n1206), .Z(n1903) );
  or2f U2044 ( .A1(n1865), .A2(n1877), .Z(n1206) );
  and2f U2054 ( .A1(n1269), .A2(n1880), .Z(n1225) );
  inv1f U2055 ( .I(n1571), .ZN(n1269) );
  or2f U2056 ( .A1(n1710), .A2(n1570), .Z(n1880) );
  or2f U2057 ( .A1(n1377), .A2(n1376), .Z(n1378) );
  or2f U2058 ( .A1(n1375), .A2(n1374), .Z(n1376) );
  or2f U2066 ( .A1(n2029), .A2(n2028), .Z(n2031) );
  and2f U2067 ( .A1(n1381), .A2(n1380), .Z(n1404) );
  and2f U2077 ( .A1(n1647), .A2(n1230), .Z(n1217) );
  or2f U2078 ( .A1(n2014), .A2(n2013), .Z(n2027) );
  and2f U2102 ( .A1(n2012), .A2(n2011), .Z(n2013) );
  or2f U2104 ( .A1(n1823), .A2(n1965), .Z(n1847) );
  and2f U2105 ( .A1(n2046), .A2(n1829), .Z(n1823) );
  or2f U2108 ( .A1(n1687), .A2(n1686), .Z(n1829) );
  and2f U2109 ( .A1(n1754), .A2(n1798), .Z(n1687) );
  and2f U2110 ( .A1(n2018), .A2(n2019), .Z(n1261) );
  and2f U2112 ( .A1(n2024), .A2(n2023), .Z(n1147) );
  or2f U2113 ( .A1(n2022), .A2(n2021), .Z(n2023) );
  or2f U2114 ( .A1(n2016), .A2(n2015), .Z(n2024) );
  or2f U2116 ( .A1(n1606), .A2(n1605), .Z(n1611) );
  or2f U2117 ( .A1(n1934), .A2(n1933), .Z(n1935) );
  and2f U2118 ( .A1(n1965), .A2(n1932), .Z(n1933) );
  or2f U2119 ( .A1(n1764), .A2(n1881), .Z(n1765) );
  and2f U2120 ( .A1(n1199), .A2(n1875), .Z(n1764) );
  or2f U2122 ( .A1(n1744), .A2(n1743), .Z(n1940) );
  and2f U2123 ( .A1(n1742), .A2(n1741), .Z(n1743) );
  inv1f U2125 ( .I(n1767), .ZN(n1864) );
  or2f U2127 ( .A1(n1182), .A2(n1183), .Z(n1767) );
  and2f U2128 ( .A1(n1270), .A2(d), .Z(n1369) );
endmodule

