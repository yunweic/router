
module too_large ( m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, 
        w, v, u, t, s, r, q, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, p0, 
        o0, n0 );
  input m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u,
         t, s, r, q, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output p0, o0, n0;
  wire   n47, n415, n421, n422, n423, n424, n425, n426, n427, n428, n429, n431,
         n432, n433, n434, n435, n436, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n494, n497, n498, n499, n500, n501, n503, n504,
         n505, n506, n507, n509, n510, n511, n513, n515, n516, n517, n518,
         n519, n520, n521, n523, n524, n525, n526, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n539, n540, n541, n542, n543,
         n544, n545, n546, n548, n549, n550, n551, n552, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025;

  or2 U30 ( .A1(u), .A2(v), .Z(n47) );
  and2 U408 ( .A1(n1025), .A2(n541), .Z(n415) );
  or2 U425 ( .A1(n536), .A2(n431), .Z(n421) );
  inv1 U426 ( .I(n764), .ZN(n422) );
  and2 U427 ( .A1(n961), .A2(n943), .Z(n423) );
  and2 U428 ( .A1(n556), .A2(n557), .Z(n424) );
  inv1 U429 ( .I(n555), .ZN(n425) );
  or2 U430 ( .A1(n785), .A2(n812), .Z(n426) );
  and2 U432 ( .A1(n999), .A2(n452), .Z(n428) );
  and2 U433 ( .A1(n511), .A2(d), .Z(n429) );
  and2 U435 ( .A1(n), .A2(o), .Z(n431) );
  or2 U436 ( .A1(n704), .A2(n520), .Z(n432) );
  and2 U440 ( .A1(n1006), .A2(n1002), .Z(n435) );
  inv1 U443 ( .I(z), .ZN(n438) );
  or2 U445 ( .A1(n924), .A2(n), .Z(n440) );
  or2 U446 ( .A1(n440), .A2(n441), .Z(n464) );
  or2 U448 ( .A1(n443), .A2(n444), .Z(n442) );
  inv1 U449 ( .I(n513), .ZN(n443) );
  inv1 U450 ( .I(n423), .ZN(n444) );
  or2 U451 ( .A1(n436), .A2(n793), .Z(n445) );
  inv1 U453 ( .I(n539), .ZN(n447) );
  or2 U455 ( .A1(n434), .A2(n802), .Z(n449) );
  or2 U456 ( .A1(n972), .A2(n924), .Z(n450) );
  inv1 U457 ( .I(n450), .ZN(n460) );
  and2 U461 ( .A1(m), .A2(b), .Z(n454) );
  inv1 U462 ( .I(n454), .ZN(n1004) );
  or2 U465 ( .A1(n525), .A2(e0), .Z(n456) );
  or2 U466 ( .A1(b0), .A2(q), .Z(n457) );
  inv1 U467 ( .I(n457), .ZN(n904) );
  and2 U470 ( .A1(o), .A2(h0), .Z(n459) );
  inv1 U471 ( .I(n459), .ZN(n562) );
  and2 U472 ( .A1(u), .A2(z), .Z(n461) );
  or2 U473 ( .A1(c0), .A2(x), .Z(n462) );
  inv1 U477 ( .I(k0), .ZN(n466) );
  and2 U478 ( .A1(n461), .A2(h0), .Z(n467) );
  and2 U480 ( .A1(m), .A2(r), .Z(n469) );
  and2 U482 ( .A1(n794), .A2(n790), .Z(n472) );
  inv1 U484 ( .I(n473), .ZN(n543) );
  inv1 U486 ( .I(n468), .ZN(n475) );
  and2 U487 ( .A1(d), .A2(k), .Z(n476) );
  inv1 U489 ( .I(n439), .ZN(n478) );
  inv1 U490 ( .I(n725), .ZN(n479) );
  or2 U494 ( .A1(n870), .A2(n546), .Z(n483) );
  and2 U495 ( .A1(n485), .A2(n657), .Z(n484) );
  inv1 U497 ( .I(n483), .ZN(n485) );
  or2 U498 ( .A1(n465), .A2(b0), .Z(n486) );
  or2 U499 ( .A1(n542), .A2(n487), .Z(n557) );
  and2 U500 ( .A1(j0), .A2(n1025), .Z(n488) );
  inv1 U501 ( .I(n488), .ZN(n487) );
  inv1 U507 ( .I(n492), .ZN(n943) );
  or2 U509 ( .A1(n818), .A2(n438), .Z(n494) );
  or2 U513 ( .A1(a0), .A2(v), .Z(n498) );
  or2 U514 ( .A1(n612), .A2(n561), .Z(n499) );
  or2 U517 ( .A1(u), .A2(n559), .Z(n501) );
  inv1 U518 ( .I(n501), .ZN(n771) );
  inv1 U521 ( .I(n934), .ZN(n504) );
  and2 U523 ( .A1(n566), .A2(n565), .Z(n506) );
  inv1 U525 ( .I(n507), .ZN(n517) );
  or2 U527 ( .A1(d0), .A2(h), .Z(n510) );
  or2 U528 ( .A1(d0), .A2(h), .Z(n509) );
  inv1 U530 ( .I(s), .ZN(n511) );
  or2 U532 ( .A1(n596), .A2(n600), .Z(n515) );
  and2 U533 ( .A1(o), .A2(h0), .Z(n516) );
  or2 U534 ( .A1(n938), .A2(j), .Z(n518) );
  and2 U537 ( .A1(n714), .A2(n713), .Z(n521) );
  or2 U538 ( .A1(n667), .A2(n668), .Z(n523) );
  and2 U543 ( .A1(n511), .A2(d), .Z(n526) );
  inv1 U544 ( .I(n429), .ZN(n973) );
  inv1 U547 ( .I(n548), .ZN(n529) );
  or2 U551 ( .A1(j0), .A2(f0), .Z(n532) );
  inv1 U552 ( .I(n532), .ZN(n580) );
  or2 U553 ( .A1(w), .A2(j), .Z(n533) );
  or2 U554 ( .A1(n920), .A2(n533), .Z(n534) );
  inv1 U555 ( .I(n534), .ZN(n994) );
  or2 U556 ( .A1(n), .A2(n562), .Z(n535) );
  inv1 U557 ( .I(n535), .ZN(n660) );
  and2 U558 ( .A1(m), .A2(r), .Z(n536) );
  inv1 U559 ( .I(n536), .ZN(n905) );
  inv1 U564 ( .I(n540), .ZN(n936) );
  inv1 U565 ( .I(y), .ZN(n541) );
  inv1 U568 ( .I(n469), .ZN(n545) );
  inv1 U569 ( .I(n545), .ZN(n546) );
  inv1 U573 ( .I(o), .ZN(n550) );
  or2 U575 ( .A1(n627), .A2(r), .Z(n551) );
  inv1 U576 ( .I(n431), .ZN(n552) );
  or2 U581 ( .A1(n1016), .A2(i0), .Z(n558) );
  inv1 U582 ( .I(d0), .ZN(n559) );
  inv1 U583 ( .I(d0), .ZN(n561) );
  inv1 U584 ( .I(d0), .ZN(n560) );
  inv1 U585 ( .I(i0), .ZN(n1025) );
  inv1 U587 ( .I(k0), .ZN(n643) );
  or2 U588 ( .A1(n643), .A2(n510), .Z(n563) );
  inv1 U589 ( .I(h0), .ZN(n793) );
  inv1 U590 ( .I(v), .ZN(n818) );
  or2 U593 ( .A1(n560), .A2(v), .Z(n564) );
  inv1 U594 ( .I(u), .ZN(n769) );
  or2 U595 ( .A1(n564), .A2(n769), .Z(n703) );
  or2 U597 ( .A1(j0), .A2(d0), .Z(n567) );
  or2 U598 ( .A1(n466), .A2(n567), .Z(n570) );
  or2 U600 ( .A1(n936), .A2(x), .Z(n568) );
  or2 U604 ( .A1(n550), .A2(d0), .Z(n571) );
  or2 U605 ( .A1(n793), .A2(n571), .Z(n572) );
  and2 U606 ( .A1(n497), .A2(n572), .Z(n573) );
  or2 U608 ( .A1(y), .A2(a0), .Z(n1016) );
  or2 U610 ( .A1(g0), .A2(f0), .Z(n577) );
  or2 U611 ( .A1(n577), .A2(e0), .Z(n961) );
  or2 U612 ( .A1(n578), .A2(n422), .Z(n610) );
  or2 U613 ( .A1(c), .A2(r), .Z(n579) );
  and2 U614 ( .A1(m), .A2(n579), .Z(n581) );
  inv1 U615 ( .I(f0), .ZN(n875) );
  inv1 U616 ( .I(h), .ZN(n845) );
  inv1 U618 ( .I(n997), .ZN(n929) );
  or2 U619 ( .A1(n581), .A2(n929), .Z(n584) );
  inv1 U620 ( .I(n), .ZN(n791) );
  or2 U621 ( .A1(n525), .A2(e0), .Z(n694) );
  or2 U622 ( .A1(n694), .A2(v), .Z(n582) );
  or2 U623 ( .A1(n582), .A2(a0), .Z(n583) );
  or2 U625 ( .A1(d0), .A2(c), .Z(n586) );
  inv1 U628 ( .I(n619), .ZN(n585) );
  or2 U629 ( .A1(n586), .A2(n585), .Z(n587) );
  or2 U630 ( .A1(n498), .A2(n561), .Z(n640) );
  or2 U632 ( .A1(n929), .A2(m), .Z(n588) );
  or2 U633 ( .A1(n588), .A2(n431), .Z(n589) );
  or2 U634 ( .A1(g), .A2(f), .Z(n590) );
  or2 U635 ( .A1(n590), .A2(e), .Z(n600) );
  or2 U638 ( .A1(n510), .A2(n1025), .Z(n593) );
  or2 U639 ( .A1(n593), .A2(c), .Z(n595) );
  or2 U640 ( .A1(n640), .A2(h), .Z(n594) );
  and2 U641 ( .A1(n595), .A2(n594), .Z(n598) );
  or2 U642 ( .A1(n596), .A2(j0), .Z(n597) );
  and2 U643 ( .A1(n598), .A2(n597), .Z(n603) );
  inv1 U645 ( .I(n925), .ZN(n796) );
  inv1 U646 ( .I(k), .ZN(n924) );
  or2 U647 ( .A1(n), .A2(n924), .Z(n971) );
  or2 U648 ( .A1(n971), .A2(n631), .Z(n599) );
  inv1 U650 ( .I(n988), .ZN(n937) );
  or2 U653 ( .A1(n601), .A2(n600), .Z(n602) );
  inv1 U656 ( .I(g0), .ZN(n607) );
  inv1 U659 ( .I(n970), .ZN(n947) );
  or2 U660 ( .A1(n491), .A2(n643), .Z(n683) );
  or2 U661 ( .A1(n608), .A2(n683), .Z(n609) );
  or2 U663 ( .A1(n562), .A2(n), .Z(n611) );
  or2 U664 ( .A1(n611), .A2(a0), .Z(n615) );
  inv1 U665 ( .I(a), .ZN(n612) );
  or2 U666 ( .A1(n499), .A2(n498), .Z(n613) );
  or2 U667 ( .A1(n613), .A2(n525), .Z(n614) );
  or2 U669 ( .A1(f0), .A2(j0), .Z(n616) );
  or2 U670 ( .A1(n616), .A2(i), .Z(n618) );
  or2 U671 ( .A1(n947), .A2(h), .Z(n617) );
  or2 U674 ( .A1(n643), .A2(d0), .Z(n620) );
  or2 U675 ( .A1(n876), .A2(n620), .Z(n621) );
  or2 U676 ( .A1(n621), .A2(n456), .Z(n622) );
  inv1 U679 ( .I(r), .ZN(n689) );
  or2 U680 ( .A1(n626), .A2(n546), .Z(n639) );
  or2 U681 ( .A1(n875), .A2(n845), .Z(n655) );
  or2 U682 ( .A1(n655), .A2(a0), .Z(n870) );
  inv1 U683 ( .I(n627), .ZN(n637) );
  and2 U684 ( .A1(k), .A2(n550), .Z(n629) );
  and2 U685 ( .A1(k), .A2(n791), .Z(n628) );
  or2 U686 ( .A1(n629), .A2(n628), .Z(n635) );
  or2 U687 ( .A1(t), .A2(l), .Z(n630) );
  inv1 U688 ( .I(n630), .ZN(n632) );
  inv1 U689 ( .I(s), .ZN(n923) );
  or2 U691 ( .A1(n632), .A2(n519), .Z(n633) );
  or2 U692 ( .A1(n633), .A2(n), .Z(n634) );
  inv1 U696 ( .I(c), .ZN(n981) );
  or2 U697 ( .A1(n640), .A2(n981), .Z(n641) );
  or2 U701 ( .A1(n763), .A2(b), .Z(n642) );
  or2 U702 ( .A1(n929), .A2(n642), .Z(n648) );
  or2 U703 ( .A1(g0), .A2(n643), .Z(n645) );
  or2 U704 ( .A1(n643), .A2(i), .Z(n644) );
  and2 U705 ( .A1(n645), .A2(n644), .Z(n646) );
  or2 U706 ( .A1(n646), .A2(n525), .Z(n647) );
  and2 U708 ( .A1(d0), .A2(a0), .Z(n649) );
  or2 U710 ( .A1(c), .A2(e), .Z(n916) );
  or2 U713 ( .A1(n650), .A2(n938), .Z(n843) );
  or2 U716 ( .A1(n654), .A2(r), .Z(n669) );
  or2 U717 ( .A1(n546), .A2(n1025), .Z(n668) );
  inv1 U718 ( .I(n655), .ZN(n656) );
  and2 U719 ( .A1(n507), .A2(n656), .Z(n658) );
  and2 U720 ( .A1(n657), .A2(n658), .Z(n666) );
  inv1 U721 ( .I(n481), .ZN(n659) );
  and2 U722 ( .A1(n552), .A2(n659), .Z(n664) );
  and2 U723 ( .A1(n550), .A2(n531), .Z(n661) );
  or2 U724 ( .A1(n661), .A2(n660), .Z(n662) );
  or2 U730 ( .A1(q), .A2(x), .Z(n673) );
  or2 U731 ( .A1(n673), .A2(b0), .Z(n941) );
  or2 U732 ( .A1(n486), .A2(y), .Z(n895) );
  and2 U734 ( .A1(n895), .A2(n675), .Z(n678) );
  and2 U735 ( .A1(n422), .A2(n895), .Z(n676) );
  or2 U736 ( .A1(n676), .A2(c0), .Z(n677) );
  inv1 U739 ( .I(n681), .ZN(n761) );
  or2 U744 ( .A1(n956), .A2(n718), .Z(n682) );
  inv1 U745 ( .I(n682), .ZN(n702) );
  inv1 U746 ( .I(n510), .ZN(n803) );
  inv1 U747 ( .I(n683), .ZN(n684) );
  and2 U748 ( .A1(n803), .A2(n684), .Z(n685) );
  and2 U749 ( .A1(n702), .A2(n685), .Z(n699) );
  or2 U751 ( .A1(n431), .A2(b), .Z(n686) );
  or2 U753 ( .A1(n525), .A2(m), .Z(n690) );
  inv1 U754 ( .I(n690), .ZN(n691) );
  and2 U756 ( .A1(n453), .A2(n693), .Z(n697) );
  or2 U757 ( .A1(n456), .A2(n546), .Z(n695) );
  inv1 U758 ( .I(n695), .ZN(n696) );
  or2 U759 ( .A1(n697), .A2(n696), .Z(n698) );
  or2 U763 ( .A1(n481), .A2(w), .Z(n711) );
  or2 U768 ( .A1(n448), .A2(n), .Z(n710) );
  or2 U772 ( .A1(n562), .A2(d0), .Z(n721) );
  inv1 U773 ( .I(x), .ZN(n907) );
  inv1 U777 ( .I(n738), .ZN(n825) );
  or2 U778 ( .A1(n825), .A2(n961), .Z(n716) );
  or2 U779 ( .A1(n716), .A2(c0), .Z(n717) );
  or2 U782 ( .A1(n469), .A2(n718), .Z(n719) );
  or2 U784 ( .A1(n734), .A2(n), .Z(n722) );
  inv1 U788 ( .I(w), .ZN(n999) );
  or2 U789 ( .A1(n561), .A2(n999), .Z(n727) );
  inv1 U790 ( .I(n727), .ZN(n740) );
  inv1 U791 ( .I(n734), .ZN(n728) );
  or2 U792 ( .A1(n480), .A2(n728), .Z(n729) );
  and2 U793 ( .A1(n552), .A2(n729), .Z(n730) );
  or2 U795 ( .A1(n455), .A2(o), .Z(n817) );
  or2 U796 ( .A1(n817), .A2(n868), .Z(n731) );
  inv1 U797 ( .I(n731), .ZN(n732) );
  or2 U800 ( .A1(n734), .A2(n768), .Z(n735) );
  or2 U801 ( .A1(n735), .A2(o), .Z(n736) );
  inv1 U802 ( .I(n736), .ZN(n754) );
  inv1 U803 ( .I(c0), .ZN(n1021) );
  inv1 U804 ( .I(n961), .ZN(n764) );
  and2 U805 ( .A1(n1021), .A2(n764), .Z(n745) );
  and2 U806 ( .A1(n415), .A2(n737), .Z(n739) );
  inv1 U808 ( .I(n768), .ZN(n741) );
  or2 U809 ( .A1(n741), .A2(n740), .Z(n742) );
  and2 U810 ( .A1(n743), .A2(n742), .Z(n744) );
  inv1 U812 ( .I(n746), .ZN(n748) );
  and2 U813 ( .A1(c), .A2(n517), .Z(n747) );
  and2 U814 ( .A1(n748), .A2(n747), .Z(n750) );
  and2 U815 ( .A1(n769), .A2(n552), .Z(n749) );
  and2 U816 ( .A1(n750), .A2(n749), .Z(n751) );
  or2 U818 ( .A1(n754), .A2(n753), .Z(n755) );
  and2 U823 ( .A1(n1021), .A2(n762), .Z(n767) );
  or2 U824 ( .A1(n467), .A2(n763), .Z(n828) );
  and2 U825 ( .A1(n764), .A2(n828), .Z(n785) );
  inv1 U826 ( .I(n486), .ZN(n765) );
  or2 U827 ( .A1(n785), .A2(n765), .Z(n766) );
  and2 U828 ( .A1(n767), .A2(n766), .Z(n784) );
  or2 U829 ( .A1(n768), .A2(n), .Z(n884) );
  or2 U830 ( .A1(n875), .A2(n845), .Z(n770) );
  and2 U833 ( .A1(h0), .A2(o), .Z(n775) );
  or2 U834 ( .A1(n775), .A2(n525), .Z(n778) );
  inv1 U835 ( .I(l0), .ZN(n848) );
  or2 U838 ( .A1(n776), .A2(i), .Z(n777) );
  and2 U840 ( .A1(n883), .A2(n885), .Z(n779) );
  or2 U844 ( .A1(n785), .A2(l0), .Z(n782) );
  and2 U847 ( .A1(n550), .A2(n545), .Z(n790) );
  inv1 U848 ( .I(j), .ZN(n989) );
  or2 U849 ( .A1(n1004), .A2(n989), .Z(n794) );
  or2 U851 ( .A1(n519), .A2(n543), .Z(n787) );
  or2 U852 ( .A1(n788), .A2(n787), .Z(n789) );
  and2 U854 ( .A1(n905), .A2(n791), .Z(n792) );
  and2 U855 ( .A1(n793), .A2(n792), .Z(n795) );
  or2 U858 ( .A1(n797), .A2(n924), .Z(n798) );
  or2 U859 ( .A1(n798), .A2(n1004), .Z(n799) );
  and2 U862 ( .A1(n803), .A2(n453), .Z(n804) );
  and2 U863 ( .A1(n490), .A2(n804), .Z(n805) );
  or2 U865 ( .A1(n546), .A2(d0), .Z(n807) );
  or2 U866 ( .A1(n), .A2(h0), .Z(n806) );
  and2 U867 ( .A1(n806), .A2(o), .Z(n874) );
  or2 U869 ( .A1(g0), .A2(n875), .Z(n808) );
  or2 U870 ( .A1(n808), .A2(e0), .Z(n809) );
  inv1 U872 ( .I(n811), .ZN(n812) );
  or2 U874 ( .A1(n455), .A2(n), .Z(n816) );
  or2 U876 ( .A1(n943), .A2(n818), .Z(n819) );
  or2 U877 ( .A1(n820), .A2(n819), .Z(n967) );
  inv1 U878 ( .I(n967), .ZN(n822) );
  or2 U881 ( .A1(n516), .A2(n825), .Z(n827) );
  or2 U882 ( .A1(n509), .A2(n848), .Z(n826) );
  or2 U883 ( .A1(n827), .A2(n826), .Z(n839) );
  inv1 U884 ( .I(n828), .ZN(n832) );
  or2 U885 ( .A1(d0), .A2(j0), .Z(n830) );
  or2 U887 ( .A1(n830), .A2(n829), .Z(n831) );
  and2 U888 ( .A1(n832), .A2(n831), .Z(n837) );
  or2 U889 ( .A1(i0), .A2(a0), .Z(n834) );
  or2 U890 ( .A1(n1025), .A2(x), .Z(n833) );
  and2 U891 ( .A1(n834), .A2(n833), .Z(n835) );
  or2 U892 ( .A1(n835), .A2(y), .Z(n836) );
  inv1 U896 ( .I(n841), .ZN(n853) );
  or2 U897 ( .A1(u), .A2(a), .Z(n842) );
  and2 U898 ( .A1(d0), .A2(n842), .Z(n844) );
  or2 U899 ( .A1(n844), .A2(n843), .Z(n850) );
  or2 U900 ( .A1(n846), .A2(n845), .Z(n847) );
  inv1 U901 ( .I(n847), .ZN(n855) );
  or2 U902 ( .A1(n855), .A2(n848), .Z(n849) );
  or2 U903 ( .A1(n850), .A2(n849), .Z(n851) );
  or2 U907 ( .A1(n855), .A2(a), .Z(n859) );
  or2 U909 ( .A1(n856), .A2(n546), .Z(n857) );
  or2 U911 ( .A1(n859), .A2(n858), .Z(n863) );
  or2 U912 ( .A1(n431), .A2(r), .Z(n861) );
  or2 U913 ( .A1(n561), .A2(n981), .Z(n860) );
  or2 U914 ( .A1(n861), .A2(n860), .Z(n862) );
  or2 U916 ( .A1(a0), .A2(u), .Z(n864) );
  or2 U917 ( .A1(n865), .A2(n864), .Z(n866) );
  or2 U919 ( .A1(n868), .A2(n), .Z(n869) );
  or2 U920 ( .A1(n869), .A2(a0), .Z(n872) );
  or2 U921 ( .A1(n870), .A2(n525), .Z(n871) );
  and2 U922 ( .A1(n872), .A2(n871), .Z(n882) );
  or2 U923 ( .A1(n874), .A2(n873), .Z(n880) );
  and2 U924 ( .A1(j0), .A2(n875), .Z(n877) );
  or2 U925 ( .A1(n877), .A2(n876), .Z(n878) );
  or2 U927 ( .A1(n878), .A2(n930), .Z(n879) );
  or2 U928 ( .A1(n880), .A2(n879), .Z(n881) );
  and2 U929 ( .A1(n882), .A2(n881), .Z(n890) );
  or2 U932 ( .A1(n886), .A2(n1025), .Z(n887) );
  and2 U937 ( .A1(n895), .A2(n894), .Z(n896) );
  or2 U938 ( .A1(n896), .A2(c0), .Z(n897) );
  and2 U943 ( .A1(n47), .A2(n492), .Z(n902) );
  inv1 U945 ( .I(n952), .ZN(n944) );
  and2 U946 ( .A1(n545), .A2(n904), .Z(n909) );
  and2 U947 ( .A1(n907), .A2(n552), .Z(n908) );
  and2 U948 ( .A1(n909), .A2(n908), .Z(n913) );
  or2 U949 ( .A1(n961), .A2(x), .Z(n910) );
  inv1 U950 ( .I(n910), .ZN(n911) );
  or2 U951 ( .A1(n911), .A2(n492), .Z(n912) );
  inv1 U954 ( .I(e0), .ZN(n1003) );
  or2 U955 ( .A1(n452), .A2(n1003), .Z(n915) );
  inv1 U956 ( .I(n915), .ZN(n940) );
  or2 U957 ( .A1(n917), .A2(n916), .Z(n918) );
  or2 U958 ( .A1(n555), .A2(n918), .Z(n919) );
  or2 U960 ( .A1(n920), .A2(j), .Z(n987) );
  and2 U962 ( .A1(k), .A2(n), .Z(n922) );
  or2 U963 ( .A1(j0), .A2(n989), .Z(n921) );
  or2 U964 ( .A1(n922), .A2(n921), .Z(n928) );
  and2 U965 ( .A1(n511), .A2(n476), .Z(n926) );
  or2 U966 ( .A1(l), .A2(t), .Z(n925) );
  inv1 U970 ( .I(m0), .ZN(n948) );
  or2 U971 ( .A1(n531), .A2(n948), .Z(n968) );
  or2 U972 ( .A1(n968), .A2(n930), .Z(n931) );
  or2 U973 ( .A1(n932), .A2(n931), .Z(n933) );
  or2 U974 ( .A1(n937), .A2(n518), .Z(n939) );
  or2 U976 ( .A1(n486), .A2(n536), .Z(n942) );
  or2 U977 ( .A1(n942), .A2(n431), .Z(n963) );
  or2 U980 ( .A1(n947), .A2(n531), .Z(n950) );
  or2 U981 ( .A1(n509), .A2(n948), .Z(n949) );
  or2 U982 ( .A1(n950), .A2(n949), .Z(n951) );
  inv1 U983 ( .I(n951), .ZN(n953) );
  or2 U984 ( .A1(n953), .A2(n952), .Z(n954) );
  inv1 U986 ( .I(n955), .ZN(n957) );
  or2 U990 ( .A1(n422), .A2(n492), .Z(n962) );
  and2 U991 ( .A1(n963), .A2(n962), .Z(n964) );
  or2 U992 ( .A1(n964), .A2(n516), .Z(n965) );
  inv1 U995 ( .I(n968), .ZN(n969) );
  and2 U996 ( .A1(n490), .A2(n969), .Z(n1012) );
  and2 U997 ( .A1(n999), .A2(n1003), .Z(n986) );
  and2 U998 ( .A1(m), .A2(n473), .Z(n975) );
  and2 U1000 ( .A1(n975), .A2(n974), .Z(n978) );
  and2 U1001 ( .A1(j), .A2(m), .Z(n976) );
  or2 U1002 ( .A1(n976), .A2(n981), .Z(n977) );
  inv1 U1005 ( .I(n980), .ZN(n998) );
  or2 U1006 ( .A1(m), .A2(n981), .Z(n982) );
  and2 U1007 ( .A1(n998), .A2(n982), .Z(n983) );
  and2 U1010 ( .A1(n989), .A2(n530), .Z(n990) );
  and2 U1012 ( .A1(n453), .A2(n425), .Z(n991) );
  or2 U1016 ( .A1(n998), .A2(n425), .Z(n1001) );
  and2 U1017 ( .A1(n428), .A2(n1001), .Z(n1008) );
  or2 U1018 ( .A1(n453), .A2(n1003), .Z(n1002) );
  or2 U1019 ( .A1(n1004), .A2(n1003), .Z(n1005) );
  and2 U1020 ( .A1(n559), .A2(n1005), .Z(n1006) );
  and2 U1021 ( .A1(n435), .A2(n1001), .Z(n1007) );
  or2 U1022 ( .A1(n1008), .A2(n1007), .Z(n1009) );
  inv1 U1027 ( .I(n1016), .ZN(n1017) );
  inv1f U424 ( .I(i), .ZN(n606) );
  inv1 U431 ( .I(j0), .ZN(n846) );
  inv1 U434 ( .I(n956), .ZN(n762) );
  or2f U437 ( .A1(n709), .A2(o), .Z(n712) );
  or2f U438 ( .A1(n715), .A2(n762), .Z(n738) );
  or2f U439 ( .A1(n607), .A2(n606), .Z(n490) );
  or2f U441 ( .A1(e0), .A2(n848), .Z(n873) );
  inv1f U442 ( .I(n531), .ZN(n868) );
  and2f U444 ( .A1(z), .A2(h0), .Z(n531) );
  or2f U447 ( .A1(i0), .A2(n846), .Z(n956) );
  or2 U452 ( .A1(n807), .A2(n874), .Z(n810) );
  or2 U454 ( .A1(n722), .A2(n721), .Z(n723) );
  and2 U458 ( .A1(n817), .A2(n816), .Z(n820) );
  or2 U459 ( .A1(n525), .A2(j), .Z(n627) );
  inv1 U460 ( .I(n773), .ZN(n763) );
  or2 U463 ( .A1(g), .A2(f), .Z(n917) );
  and2 U464 ( .A1(n618), .A2(n617), .Z(n623) );
  or2 U468 ( .A1(n874), .A2(n873), .Z(n856) );
  or2 U469 ( .A1(n516), .A2(n848), .Z(n829) );
  or2 U474 ( .A1(n1004), .A2(n796), .Z(n788) );
  or2 U475 ( .A1(n432), .A2(n433), .Z(n470) );
  and2 U476 ( .A1(n973), .A2(n468), .Z(n974) );
  and2 U479 ( .A1(w), .A2(n516), .Z(n903) );
  or2 U481 ( .A1(n491), .A2(d0), .Z(n930) );
  or2 U483 ( .A1(n584), .A2(n583), .Z(n592) );
  inv1 U485 ( .I(n484), .ZN(n638) );
  inv1 U488 ( .I(n490), .ZN(n491) );
  or2 U491 ( .A1(n752), .A2(n751), .Z(n753) );
  and2 U492 ( .A1(n888), .A2(n887), .Z(n889) );
  or2 U493 ( .A1(n883), .A2(n1025), .Z(n888) );
  and2 U496 ( .A1(n449), .A2(n805), .Z(n813) );
  or2 U502 ( .A1(n810), .A2(n809), .Z(n811) );
  or2 U503 ( .A1(n712), .A2(n711), .Z(n713) );
  or2 U504 ( .A1(n478), .A2(n479), .Z(n477) );
  or2 U505 ( .A1(n678), .A2(n677), .Z(n679) );
  inv1 U506 ( .I(n899), .ZN(n900) );
  inv1 U508 ( .I(n938), .ZN(n453) );
  and2f U510 ( .A1(n453), .A2(n1004), .Z(n452) );
  or2f U511 ( .A1(n507), .A2(n769), .Z(n481) );
  or2 U512 ( .A1(n774), .A2(n431), .Z(n883) );
  inv1 U515 ( .I(n455), .ZN(n480) );
  inv1 U516 ( .I(n549), .ZN(n505) );
  or2f U519 ( .A1(n933), .A2(n936), .Z(n549) );
  or2f U520 ( .A1(q), .A2(x), .Z(n465) );
  or2f U522 ( .A1(n528), .A2(n966), .Z(n1015) );
  or2 U524 ( .A1(n1018), .A2(n965), .Z(n966) );
  or2f U526 ( .A1(n520), .A2(n704), .Z(n463) );
  or2 U529 ( .A1(n463), .A2(n462), .Z(n706) );
  or2f U531 ( .A1(n576), .A2(n558), .Z(n556) );
  or2 U535 ( .A1(n822), .A2(n821), .Z(n823) );
  or2f U536 ( .A1(r), .A2(n462), .Z(n433) );
  or2f U539 ( .A1(n984), .A2(n983), .Z(n985) );
  or2f U540 ( .A1(n941), .A2(n421), .Z(n513) );
  or2f U541 ( .A1(n544), .A2(n551), .Z(n601) );
  inv1 U542 ( .I(n464), .ZN(n544) );
  and2f U545 ( .A1(n923), .A2(d), .Z(n631) );
  or2f U546 ( .A1(n648), .A2(n647), .Z(n651) );
  or2f U548 ( .A1(n607), .A2(n606), .Z(n970) );
  inv1 U549 ( .I(a0), .ZN(n737) );
  and2f U550 ( .A1(n587), .A2(n640), .Z(n596) );
  or2f U560 ( .A1(n901), .A2(n900), .Z(o0) );
  or2f U561 ( .A1(n824), .A2(n823), .Z(n901) );
  and2f U562 ( .A1(n795), .A2(n794), .Z(n800) );
  and2f U563 ( .A1(n791), .A2(k), .Z(n473) );
  and2f U566 ( .A1(n789), .A2(n472), .Z(n802) );
  and2f U567 ( .A1(n992), .A2(n991), .Z(n993) );
  or2f U570 ( .A1(n515), .A2(n589), .Z(n591) );
  and2f U571 ( .A1(n980), .A2(n929), .Z(n932) );
  inv1 U572 ( .I(n997), .ZN(n555) );
  inv1 U574 ( .I(n700), .ZN(n667) );
  or2f U577 ( .A1(n663), .A2(n664), .Z(n665) );
  and2f U578 ( .A1(v), .A2(n662), .Z(n663) );
  or2f U579 ( .A1(n857), .A2(n491), .Z(n858) );
  or2f U580 ( .A1(n851), .A2(n491), .Z(n852) );
  and2f U586 ( .A1(n839), .A2(n838), .Z(n840) );
  and2f U591 ( .A1(i0), .A2(n541), .Z(n540) );
  and2f U592 ( .A1(n674), .A2(n424), .Z(n675) );
  or2f U596 ( .A1(n569), .A2(n568), .Z(n674) );
  and2f U599 ( .A1(n506), .A2(n570), .Z(n569) );
  and2f U601 ( .A1(n740), .A2(n730), .Z(n733) );
  and2 U602 ( .A1(n708), .A2(n746), .Z(n448) );
  or2f U603 ( .A1(n1016), .A2(m), .Z(n707) );
  or2f U607 ( .A1(n721), .A2(n717), .Z(n724) );
  and2f U609 ( .A1(n670), .A2(n669), .Z(n524) );
  and2f U617 ( .A1(n635), .A2(n634), .Z(n636) );
  and2f U624 ( .A1(n923), .A2(d), .Z(n519) );
  or2f U626 ( .A1(l), .A2(t), .Z(n468) );
  or2f U627 ( .A1(n475), .A2(n631), .Z(n441) );
  or2f U631 ( .A1(n599), .A2(n475), .Z(n530) );
  or2f U636 ( .A1(n475), .A2(n599), .Z(n988) );
  and2f U637 ( .A1(n863), .A2(n862), .Z(n865) );
  or2f U644 ( .A1(n771), .A2(n770), .Z(n772) );
  or2f U649 ( .A1(n769), .A2(n438), .Z(n436) );
  inv1f U651 ( .I(n781), .ZN(n786) );
  and2f U652 ( .A1(n884), .A2(n779), .Z(n780) );
  or2f U654 ( .A1(n1019), .A2(n528), .Z(n1020) );
  or2f U655 ( .A1(n1018), .A2(n1017), .Z(n1019) );
  and2f U657 ( .A1(n894), .A2(n854), .Z(n867) );
  inv1 U658 ( .I(n619), .ZN(n876) );
  or2f U662 ( .A1(n649), .A2(n876), .Z(n650) );
  and2f U668 ( .A1(n425), .A2(n979), .Z(n984) );
  or2f U672 ( .A1(n978), .A2(n977), .Z(n979) );
  and2f U673 ( .A1(n708), .A2(n746), .Z(n709) );
  and2f U677 ( .A1(n521), .A2(n725), .Z(n539) );
  or2f U678 ( .A1(a0), .A2(y), .Z(n520) );
  and2f U690 ( .A1(n885), .A2(n884), .Z(n886) );
  or2f U693 ( .A1(n778), .A2(n777), .Z(n885) );
  or2f U694 ( .A1(n739), .A2(n738), .Z(n743) );
  and2f U695 ( .A1(n745), .A2(n744), .Z(n752) );
  or2f U698 ( .A1(n868), .A2(d0), .Z(n768) );
  or2f U699 ( .A1(n813), .A2(n426), .Z(n500) );
  and2f U700 ( .A1(n470), .A2(n746), .Z(n455) );
  or2f U707 ( .A1(n936), .A2(n935), .Z(n548) );
  and2f U709 ( .A1(n944), .A2(n914), .Z(n935) );
  or2f U711 ( .A1(n913), .A2(n912), .Z(n914) );
  and2f U712 ( .A1(n987), .A2(n940), .Z(n934) );
  or2f U714 ( .A1(n544), .A2(n919), .Z(n920) );
  or2f U715 ( .A1(n580), .A2(n845), .Z(n997) );
  or2f U725 ( .A1(n957), .A2(n956), .Z(n958) );
  or2f U726 ( .A1(n537), .A2(n954), .Z(n955) );
  or2f U727 ( .A1(n802), .A2(n801), .Z(n841) );
  and2f U728 ( .A1(n800), .A2(n799), .Z(n434) );
  and2f U729 ( .A1(n800), .A2(n799), .Z(n801) );
  or2f U733 ( .A1(n796), .A2(n526), .Z(n797) );
  or2f U737 ( .A1(n761), .A2(n760), .Z(n0) );
  or2f U738 ( .A1(n759), .A2(n758), .Z(n760) );
  and2f U740 ( .A1(n699), .A2(n698), .Z(n759) );
  or2f U741 ( .A1(n840), .A2(n422), .Z(n894) );
  and2f U742 ( .A1(n559), .A2(n990), .Z(n992) );
  or2f U743 ( .A1(n837), .A2(n836), .Z(n838) );
  and2f U750 ( .A1(n445), .A2(n773), .Z(n489) );
  or2f U752 ( .A1(n818), .A2(n559), .Z(n773) );
  or2f U755 ( .A1(n996), .A2(n995), .Z(n1010) );
  or2f U760 ( .A1(n993), .A2(n994), .Z(n995) );
  and2f U761 ( .A1(n986), .A2(n985), .Z(n996) );
  and2f U762 ( .A1(n940), .A2(n939), .Z(n946) );
  and2f U764 ( .A1(n945), .A2(n946), .Z(n959) );
  and2f U765 ( .A1(n442), .A2(n944), .Z(n945) );
  or2f U766 ( .A1(n916), .A2(n917), .Z(n938) );
  and2f U767 ( .A1(n605), .A2(n604), .Z(n608) );
  and2f U769 ( .A1(n592), .A2(n591), .Z(n605) );
  and2f U770 ( .A1(n565), .A2(n566), .Z(n542) );
  and2f U771 ( .A1(n563), .A2(n575), .Z(n566) );
  or2f U774 ( .A1(n559), .A2(v), .Z(n507) );
  and2f U775 ( .A1(n497), .A2(n481), .Z(n565) );
  or2f U776 ( .A1(n494), .A2(n793), .Z(n497) );
  and2f U780 ( .A1(n639), .A2(n638), .Z(n670) );
  or2f U781 ( .A1(n636), .A2(n637), .Z(n657) );
  or2f U783 ( .A1(n500), .A2(n786), .Z(n814) );
  or2f U785 ( .A1(n786), .A2(n782), .Z(n783) );
  or2f U786 ( .A1(n780), .A2(n546), .Z(n781) );
  or2f U787 ( .A1(n873), .A2(n510), .Z(n776) );
  or2f U794 ( .A1(n757), .A2(n821), .Z(n758) );
  or2f U798 ( .A1(l), .A2(t), .Z(n972) );
  and2f U799 ( .A1(n504), .A2(n505), .Z(n503) );
  or2f U807 ( .A1(n927), .A2(n928), .Z(n980) );
  or2f U811 ( .A1(n460), .A2(n926), .Z(n927) );
  or2f U817 ( .A1(n503), .A2(n529), .Z(n528) );
  or2f U819 ( .A1(n898), .A2(n897), .Z(n899) );
  or2 U820 ( .A1(n891), .A2(n546), .Z(n892) );
  and2f U821 ( .A1(n890), .A2(n889), .Z(n891) );
  and2f U822 ( .A1(n963), .A2(n423), .Z(n537) );
  inv1f U831 ( .I(n960), .ZN(n1018) );
  or2f U832 ( .A1(n959), .A2(n958), .Z(n960) );
  or2f U836 ( .A1(n902), .A2(n903), .Z(n952) );
  and2f U837 ( .A1(n999), .A2(d0), .Z(n492) );
  and2f U839 ( .A1(n1012), .A2(n1011), .Z(n1013) );
  or2f U841 ( .A1(n1010), .A2(n1009), .Z(n1011) );
  or2f U842 ( .A1(n680), .A2(n679), .Z(n681) );
  or2f U843 ( .A1(n603), .A2(n602), .Z(n604) );
  and2f U845 ( .A1(n), .A2(o), .Z(n525) );
  or2f U846 ( .A1(n692), .A2(n691), .Z(n693) );
  and2f U850 ( .A1(n689), .A2(n688), .Z(n692) );
  inv1f U853 ( .I(n458), .ZN(n688) );
  and2f U856 ( .A1(n686), .A2(n687), .Z(n458) );
  or2f U857 ( .A1(x), .A2(c0), .Z(n705) );
  or2f U860 ( .A1(n756), .A2(n755), .Z(n821) );
  or2f U861 ( .A1(n733), .A2(n732), .Z(n756) );
  or2f U864 ( .A1(n720), .A2(n719), .Z(n734) );
  and2f U868 ( .A1(n956), .A2(n936), .Z(n720) );
  or2f U871 ( .A1(n471), .A2(n705), .Z(n718) );
  or2f U873 ( .A1(q), .A2(b0), .Z(n471) );
  and2f U875 ( .A1(n1023), .A2(n1024), .Z(p0) );
  and2f U879 ( .A1(n1020), .A2(n1021), .Z(n1022) );
  and2f U880 ( .A1(n625), .A2(n624), .Z(n626) );
  and2f U886 ( .A1(n615), .A2(n614), .Z(n625) );
  or2f U893 ( .A1(n623), .A2(n622), .Z(n624) );
  and2f U894 ( .A1(n672), .A2(n671), .Z(n680) );
  and2f U895 ( .A1(n524), .A2(n523), .Z(n671) );
  and2f U904 ( .A1(n610), .A2(n609), .Z(n672) );
  or2f U905 ( .A1(n726), .A2(n477), .Z(n757) );
  and2f U906 ( .A1(n702), .A2(n701), .Z(n726) );
  and2f U908 ( .A1(n700), .A2(n545), .Z(n701) );
  or2f U910 ( .A1(n666), .A2(n665), .Z(n700) );
  or2f U915 ( .A1(n853), .A2(n852), .Z(n854) );
  and2f U918 ( .A1(n893), .A2(n892), .Z(n898) );
  and2f U926 ( .A1(n867), .A2(n866), .Z(n893) );
  or2f U930 ( .A1(i0), .A2(n737), .Z(n619) );
  and2f U931 ( .A1(n815), .A2(n814), .Z(n824) );
  and2f U933 ( .A1(n783), .A2(n784), .Z(n815) );
  and2f U934 ( .A1(n489), .A2(n772), .Z(n774) );
  or2f U935 ( .A1(n706), .A2(r), .Z(n708) );
  or2f U936 ( .A1(n707), .A2(n718), .Z(n746) );
  and2f U939 ( .A1(n714), .A2(n713), .Z(n439) );
  or2f U940 ( .A1(n711), .A2(n710), .Z(n714) );
  or2f U941 ( .A1(q), .A2(b0), .Z(n704) );
  or2f U942 ( .A1(n1014), .A2(n1015), .Z(n1024) );
  or2f U944 ( .A1(n1013), .A2(n446), .Z(n1014) );
  or2f U952 ( .A1(n1022), .A2(n446), .Z(n1023) );
  or2f U953 ( .A1(n447), .A2(n822), .Z(n446) );
  and2f U959 ( .A1(n907), .A2(n540), .Z(n715) );
  and2f U961 ( .A1(n724), .A2(n723), .Z(n725) );
  and2f U967 ( .A1(n653), .A2(n652), .Z(n654) );
  or2f U968 ( .A1(n641), .A2(n687), .Z(n653) );
  or2f U969 ( .A1(n651), .A2(n843), .Z(n652) );
  or2f U975 ( .A1(n544), .A2(n627), .Z(n687) );
  and2f U978 ( .A1(n703), .A2(n570), .Z(n574) );
  and2f U979 ( .A1(n574), .A2(n575), .Z(n482) );
  or2f U985 ( .A1(n562), .A2(n818), .Z(n575) );
  and2f U987 ( .A1(n482), .A2(n573), .Z(n576) );
  and2f U988 ( .A1(n427), .A2(n674), .Z(n578) );
  and2f U989 ( .A1(n556), .A2(n557), .Z(n427) );
endmodule

