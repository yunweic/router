
module C499_iscas ( o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, 
        z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, 
        b, a, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, 
        e1, d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0 );
  input o0, n0, m0, l0, k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w,
         v, u, t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1,
         d1, c1, b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0;
  wire   n499, n500, n501, n502, n503, n505, n506, n507, n508, n509, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n533, n534, n535,
         n537, n538, n539, n540, n541, n542, n543, n545, n546, n548, n549,
         n550, n551, n553, n554, n555, n556, n558, n561, n562, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n632, n633, n634,
         n635, n637, n638, n639, n641, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n656, n657, n658, n659, n661,
         n662, n663, n664, n665, n666, n667, n670, n671, n674, n675, n676,
         n677, n678, n680, n681, n683, n684, n685, n686, n687, n688, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1033,
         n1034, n1035, n1036, n1037, n1038, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1073, n1074, n1075,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1086, n1087,
         n1088, n1089, n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1126, n1127, n1128, n1129, n1130,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197;

  or2 U537 ( .A1(n499), .A2(n624), .Z(n505) );
  inv1 U546 ( .I(n624), .ZN(n514) );
  inv1 U547 ( .I(n514), .ZN(n515) );
  and2 U557 ( .A1(n724), .A2(n723), .Z(n525) );
  and2 U561 ( .A1(n930), .A2(n531), .Z(n529) );
  and2 U567 ( .A1(n753), .A2(n667), .Z(n534) );
  or2 U570 ( .A1(n720), .A2(n723), .Z(n537) );
  inv1 U575 ( .I(n1158), .ZN(n541) );
  inv1 U579 ( .I(n888), .ZN(n545) );
  or2 U585 ( .A1(n512), .A2(n818), .Z(n550) );
  or2 U590 ( .A1(n727), .A2(n730), .Z(n555) );
  inv1 U606 ( .I(n895), .ZN(n568) );
  inv1 U612 ( .I(e), .ZN(n573) );
  inv1 U619 ( .I(n599), .ZN(n580) );
  inv1 U620 ( .I(c0), .ZN(n581) );
  or2 U623 ( .A1(n586), .A2(n648), .Z(n584) );
  inv1 U630 ( .I(n588), .ZN(n890) );
  inv1 U633 ( .I(o), .ZN(n590) );
  inv1 U635 ( .I(f), .ZN(n592) );
  or2 U639 ( .A1(n795), .A2(n798), .Z(n596) );
  or2 U641 ( .A1(n1195), .A2(n598), .Z(n1173) );
  or2 U642 ( .A1(n542), .A2(n685), .Z(n598) );
  or2 U658 ( .A1(n902), .A2(n578), .Z(n615) );
  or2 U659 ( .A1(n953), .A2(n617), .Z(n616) );
  inv1 U661 ( .I(n954), .ZN(n617) );
  inv1 U664 ( .I(r), .ZN(n619) );
  and2 U667 ( .A1(n930), .A2(n929), .Z(n622) );
  inv1 U672 ( .I(n625), .ZN(n961) );
  inv1 U676 ( .I(n759), .ZN(n628) );
  inv1 U697 ( .I(n647), .ZN(n664) );
  inv1 U698 ( .I(n1129), .ZN(n648) );
  inv1 U699 ( .I(v), .ZN(n649) );
  or2 U700 ( .A1(n767), .A2(n766), .Z(n650) );
  inv1 U703 ( .I(h), .ZN(n653) );
  inv1 U705 ( .I(n654), .ZN(n686) );
  or2 U709 ( .A1(n579), .A2(n865), .Z(n657) );
  or2 U714 ( .A1(n863), .A2(n663), .Z(n662) );
  inv1 U716 ( .I(n864), .ZN(n663) );
  inv1 U718 ( .I(n665), .ZN(n794) );
  inv1 U719 ( .I(n793), .ZN(n666) );
  or2 U731 ( .A1(n644), .A2(n1124), .Z(n678) );
  inv1 U738 ( .I(p), .ZN(n687) );
  and2 U742 ( .A1(o), .A2(n620), .Z(n691) );
  inv1 U743 ( .I(o), .ZN(n1059) );
  and2 U744 ( .A1(n1059), .A2(k), .Z(n690) );
  or2 U745 ( .A1(n691), .A2(n690), .Z(n695) );
  inv1 U746 ( .I(c), .ZN(n976) );
  and2 U747 ( .A1(g), .A2(n976), .Z(n693) );
  and2 U749 ( .A1(n1004), .A2(c), .Z(n692) );
  or2 U750 ( .A1(n693), .A2(n692), .Z(n696) );
  inv1 U751 ( .I(n696), .ZN(n694) );
  and2 U752 ( .A1(n695), .A2(n694), .Z(n699) );
  inv1 U753 ( .I(n695), .ZN(n697) );
  and2 U754 ( .A1(n697), .A2(n696), .Z(n698) );
  or2 U755 ( .A1(n699), .A2(n698), .Z(n728) );
  inv1 U758 ( .I(t), .ZN(n1097) );
  inv1 U761 ( .I(q), .ZN(n1079) );
  inv1 U771 ( .I(n754), .ZN(n753) );
  inv1 U772 ( .I(a0), .ZN(n1147) );
  inv1 U777 ( .I(y), .ZN(n1135) );
  inv1 U791 ( .I(o0), .ZN(n952) );
  inv1 U792 ( .I(i0), .ZN(n722) );
  or2 U793 ( .A1(n952), .A2(n722), .Z(n725) );
  inv1 U794 ( .I(n725), .ZN(n723) );
  inv1 U797 ( .I(n728), .ZN(n730) );
  and2 U800 ( .A1(n1020), .A2(m), .Z(n734) );
  inv1 U801 ( .I(m), .ZN(n1047) );
  and2 U802 ( .A1(i), .A2(n1047), .Z(n733) );
  or2 U803 ( .A1(n734), .A2(n733), .Z(n738) );
  inv1 U804 ( .I(a), .ZN(n964) );
  and2 U805 ( .A1(e), .A2(n964), .Z(n736) );
  inv1 U806 ( .I(e), .ZN(n992) );
  and2 U807 ( .A1(n992), .A2(a), .Z(n735) );
  or2 U808 ( .A1(n736), .A2(n735), .Z(n739) );
  inv1 U809 ( .I(n739), .ZN(n737) );
  and2 U810 ( .A1(n738), .A2(n737), .Z(n742) );
  inv1 U811 ( .I(n738), .ZN(n740) );
  and2 U812 ( .A1(n740), .A2(n739), .Z(n741) );
  or2 U813 ( .A1(n742), .A2(n741), .Z(n763) );
  inv1 U814 ( .I(w), .ZN(n1119) );
  inv1 U819 ( .I(u), .ZN(n1107) );
  inv1 U821 ( .I(v), .ZN(n1113) );
  inv1 U833 ( .I(g0), .ZN(n757) );
  or2 U834 ( .A1(n757), .A2(n952), .Z(n759) );
  inv1 U839 ( .I(n763), .ZN(n765) );
  inv1 U845 ( .I(n), .ZN(n1053) );
  and2 U846 ( .A1(n1053), .A2(j), .Z(n768) );
  or2 U847 ( .A1(n769), .A2(n768), .Z(n773) );
  and2 U849 ( .A1(f), .A2(n570), .Z(n771) );
  inv1 U850 ( .I(f), .ZN(n998) );
  and2 U851 ( .A1(n998), .A2(b), .Z(n770) );
  or2 U852 ( .A1(n771), .A2(n770), .Z(n774) );
  inv1 U853 ( .I(n774), .ZN(n772) );
  and2 U854 ( .A1(n773), .A2(n772), .Z(n777) );
  inv1 U855 ( .I(n773), .ZN(n775) );
  and2 U856 ( .A1(n775), .A2(n774), .Z(n776) );
  or2 U857 ( .A1(n777), .A2(n776), .Z(n796) );
  inv1 U858 ( .I(e0), .ZN(n1174) );
  inv1 U859 ( .I(f0), .ZN(n1181) );
  inv1 U862 ( .I(c0), .ZN(n1162) );
  inv1 U864 ( .I(d0), .ZN(n1169) );
  and2 U865 ( .A1(n633), .A2(c0), .Z(n779) );
  inv1 U876 ( .I(h0), .ZN(n791) );
  or2 U877 ( .A1(n952), .A2(n791), .Z(n793) );
  inv1 U880 ( .I(n796), .ZN(n798) );
  and2 U884 ( .A1(p), .A2(n614), .Z(n802) );
  inv1 U885 ( .I(p), .ZN(n1067) );
  and2 U886 ( .A1(n1067), .A2(l), .Z(n801) );
  or2 U887 ( .A1(n802), .A2(n801), .Z(n806) );
  and2 U889 ( .A1(h), .A2(n605), .Z(n804) );
  inv1 U890 ( .I(h), .ZN(n1011) );
  and2 U891 ( .A1(n1011), .A2(d), .Z(n803) );
  or2 U892 ( .A1(n804), .A2(n803), .Z(n807) );
  inv1 U893 ( .I(n807), .ZN(n805) );
  and2 U894 ( .A1(n806), .A2(n805), .Z(n810) );
  inv1 U895 ( .I(n806), .ZN(n808) );
  and2 U896 ( .A1(n808), .A2(n807), .Z(n809) );
  or2 U897 ( .A1(n810), .A2(n809), .Z(n823) );
  inv1 U901 ( .I(j0), .ZN(n817) );
  or2 U902 ( .A1(n952), .A2(n817), .Z(n820) );
  inv1 U903 ( .I(n820), .ZN(n818) );
  inv1 U906 ( .I(n823), .ZN(n825) );
  and2 U915 ( .A1(n1154), .A2(f0), .Z(n832) );
  and2 U916 ( .A1(b0), .A2(n1181), .Z(n831) );
  or2 U917 ( .A1(n832), .A2(n831), .Z(n836) );
  and2 U918 ( .A1(n1097), .A2(x), .Z(n834) );
  and2 U919 ( .A1(t), .A2(n600), .Z(n833) );
  or2 U920 ( .A1(n834), .A2(n833), .Z(n837) );
  inv1 U921 ( .I(n837), .ZN(n835) );
  and2 U922 ( .A1(n836), .A2(n835), .Z(n840) );
  inv1 U923 ( .I(n836), .ZN(n838) );
  and2 U924 ( .A1(n838), .A2(n837), .Z(n839) );
  or2 U925 ( .A1(n840), .A2(n839), .Z(n867) );
  inv1 U951 ( .I(n0), .ZN(n862) );
  or2 U952 ( .A1(n952), .A2(n862), .Z(n864) );
  inv1 U955 ( .I(n867), .ZN(n869) );
  and2 U959 ( .A1(n645), .A2(d0), .Z(n873) );
  and2 U960 ( .A1(z), .A2(n1169), .Z(n872) );
  or2 U961 ( .A1(n873), .A2(n872), .Z(n877) );
  and2 U962 ( .A1(n619), .A2(v), .Z(n875) );
  and2 U963 ( .A1(r), .A2(n1113), .Z(n874) );
  or2 U964 ( .A1(n875), .A2(n874), .Z(n878) );
  inv1 U965 ( .I(n878), .ZN(n876) );
  and2 U966 ( .A1(n877), .A2(n876), .Z(n881) );
  inv1 U967 ( .I(n877), .ZN(n879) );
  and2 U968 ( .A1(n879), .A2(n878), .Z(n880) );
  or2 U969 ( .A1(n881), .A2(n880), .Z(n899) );
  inv1 U970 ( .I(l0), .ZN(n882) );
  or2 U971 ( .A1(n952), .A2(n882), .Z(n895) );
  or2 U977 ( .A1(n886), .A2(n885), .Z(n888) );
  inv1 U984 ( .I(n899), .ZN(n901) );
  and2 U988 ( .A1(n1135), .A2(c0), .Z(n904) );
  and2 U989 ( .A1(y), .A2(n1162), .Z(n903) );
  or2 U990 ( .A1(n904), .A2(n903), .Z(n908) );
  and2 U991 ( .A1(n1079), .A2(u), .Z(n906) );
  and2 U992 ( .A1(q), .A2(n1107), .Z(n905) );
  or2 U993 ( .A1(n906), .A2(n905), .Z(n909) );
  inv1 U994 ( .I(n909), .ZN(n907) );
  and2 U995 ( .A1(n908), .A2(n907), .Z(n912) );
  and2 U997 ( .A1(n910), .A2(n909), .Z(n911) );
  or2 U998 ( .A1(n912), .A2(n911), .Z(n933) );
  inv1 U1014 ( .I(k0), .ZN(n926) );
  or2 U1015 ( .A1(n952), .A2(n926), .Z(n929) );
  inv1 U1016 ( .I(n929), .ZN(n927) );
  inv1 U1021 ( .I(n933), .ZN(n935) );
  and2 U1024 ( .A1(n1147), .A2(e0), .Z(n938) );
  and2 U1025 ( .A1(a0), .A2(n1174), .Z(n937) );
  or2 U1026 ( .A1(n938), .A2(n937), .Z(n942) );
  and2 U1027 ( .A1(n612), .A2(w), .Z(n940) );
  and2 U1028 ( .A1(s), .A2(n1119), .Z(n939) );
  or2 U1029 ( .A1(n940), .A2(n939), .Z(n943) );
  inv1 U1030 ( .I(n943), .ZN(n941) );
  and2 U1031 ( .A1(n942), .A2(n941), .Z(n946) );
  inv1 U1032 ( .I(n942), .ZN(n944) );
  and2 U1033 ( .A1(n944), .A2(n943), .Z(n945) );
  or2 U1034 ( .A1(n946), .A2(n945), .Z(n957) );
  inv1 U1038 ( .I(m0), .ZN(n951) );
  or2 U1039 ( .A1(n952), .A2(n951), .Z(n954) );
  inv1 U1042 ( .I(n957), .ZN(n959) );
  or2 U1045 ( .A1(n980), .A2(n586), .Z(n962) );
  or2 U1048 ( .A1(n963), .A2(a), .Z(n967) );
  and2 U1050 ( .A1(n967), .A2(n966), .Z(p0) );
  or2 U1051 ( .A1(n626), .A2(n520), .Z(n968) );
  or2 U1054 ( .A1(n969), .A2(b), .Z(n973) );
  and2 U1056 ( .A1(n973), .A2(n972), .Z(q0) );
  or2 U1057 ( .A1(n980), .A2(n1194), .Z(n974) );
  inv1 U1059 ( .I(n977), .ZN(n975) );
  or2 U1060 ( .A1(n975), .A2(c), .Z(n979) );
  or2 U1061 ( .A1(n977), .A2(n976), .Z(n978) );
  and2 U1062 ( .A1(n979), .A2(n978), .Z(r0) );
  inv1 U1065 ( .I(n984), .ZN(n982) );
  or2 U1066 ( .A1(n982), .A2(d), .Z(n986) );
  or2 U1067 ( .A1(n984), .A2(n605), .Z(n985) );
  and2 U1068 ( .A1(n986), .A2(n985), .Z(s0) );
  or2 U1077 ( .A1(n993), .A2(n992), .Z(n994) );
  and2 U1078 ( .A1(n995), .A2(n994), .Z(t0) );
  or2 U1079 ( .A1(n1008), .A2(n520), .Z(n996) );
  or2 U1082 ( .A1(n997), .A2(f), .Z(n1001) );
  and2 U1084 ( .A1(n1001), .A2(n1000), .Z(u0) );
  or2 U1085 ( .A1(n516), .A2(n1194), .Z(n1002) );
  inv1 U1087 ( .I(n1005), .ZN(n1003) );
  or2 U1088 ( .A1(n1003), .A2(g), .Z(n1007) );
  or2 U1089 ( .A1(n1005), .A2(n1004), .Z(n1006) );
  and2 U1090 ( .A1(n1007), .A2(n1006), .Z(v0) );
  inv1 U1093 ( .I(n1012), .ZN(n1010) );
  or2 U1094 ( .A1(n1010), .A2(h), .Z(n1014) );
  or2 U1095 ( .A1(n1012), .A2(n1011), .Z(n1013) );
  and2 U1096 ( .A1(n1014), .A2(n1013), .Z(w0) );
  or2 U1101 ( .A1(n594), .A2(n586), .Z(n1018) );
  or2 U1104 ( .A1(n1019), .A2(i), .Z(n1023) );
  or2 U1105 ( .A1(n1021), .A2(n1020), .Z(n1022) );
  and2 U1106 ( .A1(n1023), .A2(n1022), .Z(x0) );
  or2 U1110 ( .A1(n1025), .A2(j), .Z(n1029) );
  or2 U1111 ( .A1(n1027), .A2(n1026), .Z(n1028) );
  and2 U1112 ( .A1(n1029), .A2(n1028), .Z(y0) );
  or2 U1113 ( .A1(n1036), .A2(n1194), .Z(n1030) );
  or2 U1116 ( .A1(n1031), .A2(k), .Z(n1035) );
  or2 U1117 ( .A1(n1033), .A2(n620), .Z(n1034) );
  and2 U1118 ( .A1(n1035), .A2(n1034), .Z(z0) );
  or2 U1119 ( .A1(n594), .A2(n648), .Z(n1037) );
  or2 U1123 ( .A1(n1040), .A2(n614), .Z(n1041) );
  and2 U1124 ( .A1(n1042), .A2(n1041), .Z(a1) );
  or2 U1127 ( .A1(n1063), .A2(n586), .Z(n1045) );
  or2 U1130 ( .A1(n1046), .A2(m), .Z(n1050) );
  or2 U1131 ( .A1(n1048), .A2(n1047), .Z(n1049) );
  and2 U1132 ( .A1(n1050), .A2(n1049), .Z(b1) );
  or2 U1133 ( .A1(n1063), .A2(n520), .Z(n1051) );
  or2 U1136 ( .A1(n1052), .A2(n), .Z(n1056) );
  or2 U1137 ( .A1(n1054), .A2(n1053), .Z(n1055) );
  and2 U1138 ( .A1(n1056), .A2(n1055), .Z(c1) );
  inv1 U1141 ( .I(n1060), .ZN(n1058) );
  or2 U1142 ( .A1(n1058), .A2(o), .Z(n1062) );
  or2 U1143 ( .A1(n1060), .A2(n1059), .Z(n1061) );
  and2 U1144 ( .A1(n1062), .A2(n1061), .Z(d1) );
  or2 U1145 ( .A1(n513), .A2(n648), .Z(n1065) );
  or2 U1148 ( .A1(n1066), .A2(p), .Z(n1070) );
  or2 U1149 ( .A1(n1068), .A2(n1067), .Z(n1069) );
  and2 U1150 ( .A1(n1070), .A2(n1069), .Z(e1) );
  or2 U1157 ( .A1(n1078), .A2(q), .Z(n1082) );
  or2 U1158 ( .A1(n1080), .A2(n1079), .Z(n1081) );
  and2 U1159 ( .A1(n1082), .A2(n1081), .Z(f1) );
  or2 U1163 ( .A1(n1084), .A2(r), .Z(n1088) );
  or2 U1164 ( .A1(n1086), .A2(n619), .Z(n1087) );
  and2 U1165 ( .A1(n1088), .A2(n1087), .Z(g1) );
  or2 U1169 ( .A1(n1090), .A2(s), .Z(n1094) );
  or2 U1170 ( .A1(n612), .A2(n1092), .Z(n1093) );
  and2 U1171 ( .A1(n1094), .A2(n1093), .Z(h1) );
  or2 U1175 ( .A1(n1096), .A2(t), .Z(n1100) );
  or2 U1176 ( .A1(n1098), .A2(n1097), .Z(n1099) );
  and2 U1177 ( .A1(n1100), .A2(n1099), .Z(i1) );
  inv1 U1181 ( .I(n1108), .ZN(n1106) );
  or2 U1182 ( .A1(n1106), .A2(u), .Z(n1110) );
  or2 U1183 ( .A1(n1108), .A2(n1107), .Z(n1109) );
  and2 U1184 ( .A1(n1110), .A2(n1109), .Z(j1) );
  inv1 U1187 ( .I(n1114), .ZN(n1112) );
  or2 U1188 ( .A1(n1112), .A2(v), .Z(n1116) );
  or2 U1189 ( .A1(n1114), .A2(n1113), .Z(n1115) );
  and2 U1190 ( .A1(n1116), .A2(n1115), .Z(k1) );
  or2 U1194 ( .A1(n1118), .A2(w), .Z(n1122) );
  or2 U1195 ( .A1(n1120), .A2(n1119), .Z(n1121) );
  and2 U1196 ( .A1(n1122), .A2(n1121), .Z(l1) );
  or2 U1199 ( .A1(n664), .A2(x), .Z(n1126) );
  and2 U1200 ( .A1(n1126), .A2(n1127), .Z(m1) );
  inv1 U1205 ( .I(n1136), .ZN(n1134) );
  or2 U1206 ( .A1(n1134), .A2(y), .Z(n1138) );
  or2 U1207 ( .A1(n1136), .A2(n1135), .Z(n1137) );
  and2 U1208 ( .A1(n1138), .A2(n1137), .Z(n1) );
  or2 U1212 ( .A1(n1140), .A2(z), .Z(n1144) );
  and2 U1214 ( .A1(n1144), .A2(n1143), .Z(o1) );
  or2 U1215 ( .A1(n1151), .A2(n685), .Z(n1145) );
  or2 U1219 ( .A1(n1148), .A2(n1147), .Z(n1149) );
  and2 U1220 ( .A1(n1150), .A2(n1149), .Z(p1) );
  or2 U1224 ( .A1(n1153), .A2(b0), .Z(n1157) );
  or2 U1225 ( .A1(n1155), .A2(n1154), .Z(n1156) );
  and2 U1226 ( .A1(n1157), .A2(n1156), .Z(q1) );
  or2 U1230 ( .A1(n1161), .A2(c0), .Z(n1165) );
  or2 U1231 ( .A1(n1163), .A2(n1162), .Z(n1164) );
  and2 U1232 ( .A1(n1165), .A2(n1164), .Z(r1) );
  or2 U1236 ( .A1(n1168), .A2(d0), .Z(n1172) );
  or2 U1237 ( .A1(n1170), .A2(n1169), .Z(n1171) );
  and2 U1238 ( .A1(n1172), .A2(n1171), .Z(s1) );
  or2 U1240 ( .A1(n654), .A2(n1174), .Z(n1175) );
  and2 U1241 ( .A1(n1176), .A2(n1175), .Z(t1) );
  or2 U1245 ( .A1(n1180), .A2(f0), .Z(n1184) );
  or2 U1246 ( .A1(n1182), .A2(n1181), .Z(n1183) );
  and2 U1247 ( .A1(n1184), .A2(n1183), .Z(u1) );
  inv1 U653 ( .I(n561), .ZN(n1185) );
  inv1f U530 ( .I(s), .ZN(n612) );
  inv1f U531 ( .I(n548), .ZN(n602) );
  inv1f U532 ( .I(b0), .ZN(n1154) );
  inv1f U533 ( .I(n602), .ZN(n586) );
  inv1f U534 ( .I(z), .ZN(n645) );
  inv1 U535 ( .I(n), .ZN(n643) );
  inv1 U536 ( .I(m), .ZN(n593) );
  and2 U538 ( .A1(n597), .A2(v), .Z(n521) );
  inv1 U539 ( .I(n782), .ZN(n784) );
  inv1 U540 ( .I(n567), .ZN(n898) );
  inv1 U541 ( .I(n630), .ZN(n1129) );
  inv1 U542 ( .I(n675), .ZN(n827) );
  or2f U543 ( .A1(n816), .A2(n815), .Z(n819) );
  and2 U544 ( .A1(n819), .A2(n818), .Z(n571) );
  or2f U545 ( .A1(n827), .A2(n826), .Z(n1102) );
  inv1f U548 ( .I(n1080), .ZN(n1078) );
  inv1f U549 ( .I(n1155), .ZN(n1153) );
  inv1f U550 ( .I(n1182), .ZN(n1180) );
  and2f U551 ( .A1(d0), .A2(n581), .Z(n780) );
  or2f U552 ( .A1(n752), .A2(n528), .Z(n637) );
  and2f U553 ( .A1(n1189), .A2(n566), .Z(n1192) );
  and2f U554 ( .A1(n824), .A2(n825), .Z(n522) );
  or2f U555 ( .A1(n711), .A2(n710), .Z(n715) );
  inv1f U556 ( .I(n540), .ZN(n1193) );
  inv1 U558 ( .I(n928), .ZN(n930) );
  or2 U559 ( .A1(n516), .A2(n586), .Z(n990) );
  inv1 U560 ( .I(n846), .ZN(n844) );
  inv1 U562 ( .I(n845), .ZN(n847) );
  inv1 U563 ( .I(n856), .ZN(n854) );
  inv1 U564 ( .I(n715), .ZN(n717) );
  or2 U565 ( .A1(n713), .A2(n712), .Z(n517) );
  inv1 U566 ( .I(n748), .ZN(n750) );
  or2 U568 ( .A1(n521), .A2(n745), .Z(n572) );
  inv1 U569 ( .I(n783), .ZN(n781) );
  inv1 U571 ( .I(n749), .ZN(n747) );
  and2 U572 ( .A1(n597), .A2(v), .Z(n746) );
  and2 U573 ( .A1(n889), .A2(n527), .Z(n549) );
  and2 U574 ( .A1(n), .A2(n1026), .Z(n769) );
  inv1 U576 ( .I(n908), .ZN(n910) );
  inv1 U577 ( .I(n606), .ZN(n987) );
  inv1 U578 ( .I(n658), .ZN(n508) );
  or2 U580 ( .A1(n632), .A2(n548), .Z(n499) );
  or2 U581 ( .A1(n630), .A2(n548), .Z(n1103) );
  and2 U582 ( .A1(n900), .A2(n901), .Z(n1186) );
  inv1 U583 ( .I(d), .ZN(n605) );
  or2 U584 ( .A1(n1008), .A2(n648), .Z(n1009) );
  or2 U586 ( .A1(n1036), .A2(n520), .Z(n1024) );
  inv1 U587 ( .I(x), .ZN(n600) );
  or2 U588 ( .A1(n991), .A2(e), .Z(n995) );
  or2 U589 ( .A1(n1038), .A2(l), .Z(n1042) );
  inv1 U591 ( .I(n1086), .ZN(n1084) );
  inv1 U592 ( .I(n1098), .ZN(n1096) );
  inv1 U593 ( .I(n1120), .ZN(n1118) );
  or2 U594 ( .A1(n1142), .A2(n645), .Z(n1143) );
  inv1 U595 ( .I(n1148), .ZN(n1146) );
  inv1 U596 ( .I(n1163), .ZN(n1161) );
  inv1 U597 ( .I(n1170), .ZN(n1168) );
  or2 U598 ( .A1(n686), .A2(e0), .Z(n1176) );
  inv1 U599 ( .I(n676), .ZN(n1194) );
  inv1 U600 ( .I(n656), .ZN(n676) );
  or2 U601 ( .A1(n932), .A2(n935), .Z(n623) );
  and2f U602 ( .A1(n507), .A2(n927), .Z(n932) );
  inv1f U603 ( .I(l), .ZN(n614) );
  or2f U604 ( .A1(n1128), .A2(n641), .Z(n1195) );
  inv1f U605 ( .I(k), .ZN(n620) );
  and2f U607 ( .A1(n830), .A2(n829), .Z(n1196) );
  or2 U608 ( .A1(n971), .A2(n570), .Z(n972) );
  or2 U609 ( .A1(n965), .A2(n964), .Z(n966) );
  and2f U610 ( .A1(n830), .A2(n564), .Z(n1197) );
  or2 U611 ( .A1(n999), .A2(n998), .Z(n1000) );
  inv1f U613 ( .I(n538), .ZN(n1044) );
  inv1f U614 ( .I(n1071), .ZN(n1188) );
  inv1f U615 ( .I(n1142), .ZN(n1140) );
  inv1f U616 ( .I(n971), .ZN(n969) );
  inv1f U617 ( .I(n965), .ZN(n963) );
  inv1f U618 ( .I(n1027), .ZN(n1025) );
  inv1f U621 ( .I(n999), .ZN(n997) );
  inv1f U622 ( .I(n587), .ZN(n732) );
  inv1f U624 ( .I(n632), .ZN(n641) );
  or2f U625 ( .A1(n1104), .A2(n515), .Z(n585) );
  inv1 U626 ( .I(b), .ZN(n570) );
  or2 U627 ( .A1(n709), .A2(n708), .Z(n674) );
  inv1 U628 ( .I(n887), .ZN(n889) );
  or2f U629 ( .A1(n866), .A2(n869), .Z(n579) );
  and2 U631 ( .A1(n863), .A2(n663), .Z(n866) );
  or2f U632 ( .A1(n555), .A2(n726), .Z(n587) );
  or2f U634 ( .A1(n1104), .A2(n1103), .Z(n1123) );
  inv1f U636 ( .I(n813), .ZN(n811) );
  inv1f U637 ( .I(d0), .ZN(n633) );
  or2f U638 ( .A1(n865), .A2(n866), .Z(n868) );
  inv1 U640 ( .I(n662), .ZN(n865) );
  and2f U643 ( .A1(n857), .A2(n562), .Z(n577) );
  inv1f U644 ( .I(n1033), .ZN(n1031) );
  inv1f U645 ( .I(n1048), .ZN(n1046) );
  or2f U646 ( .A1(n752), .A2(n528), .Z(n812) );
  or2f U647 ( .A1(n902), .A2(n535), .Z(n606) );
  and2f U648 ( .A1(k), .A2(n614), .Z(n884) );
  and2f U649 ( .A1(n1154), .A2(a0), .Z(n710) );
  and2f U650 ( .A1(n762), .A2(n763), .Z(n638) );
  inv1f U651 ( .I(n1187), .ZN(n762) );
  and2f U652 ( .A1(n762), .A2(n763), .Z(n767) );
  inv1f U654 ( .I(n657), .ZN(n871) );
  or2f U655 ( .A1(n859), .A2(n577), .Z(n688) );
  inv1f U656 ( .I(n677), .ZN(n821) );
  and2f U657 ( .A1(n620), .A2(l), .Z(n883) );
  inv1f U660 ( .I(n616), .ZN(n955) );
  or2f U662 ( .A1(n595), .A2(n955), .Z(n625) );
  and2f U663 ( .A1(n958), .A2(n959), .Z(n960) );
  inv1f U665 ( .I(n1092), .ZN(n1090) );
  or2f U666 ( .A1(n956), .A2(n959), .Z(n595) );
  or2f U668 ( .A1(n613), .A2(n1166), .Z(n1167) );
  and2f U669 ( .A1(n901), .A2(n900), .Z(n578) );
  or2f U670 ( .A1(n613), .A2(n515), .Z(n1160) );
  inv1f U671 ( .I(n1054), .ZN(n1052) );
  and2 U673 ( .A1(n935), .A2(n934), .Z(n609) );
  and2 U674 ( .A1(n934), .A2(n935), .Z(n936) );
  and2 U675 ( .A1(n935), .A2(n533), .Z(n530) );
  and2f U677 ( .A1(n929), .A2(n935), .Z(n531) );
  and2f U678 ( .A1(b0), .A2(n1147), .Z(n711) );
  or2f U679 ( .A1(n732), .A2(n731), .Z(n656) );
  and2f U680 ( .A1(n729), .A2(n730), .Z(n731) );
  or2f U681 ( .A1(n600), .A2(n678), .Z(n1127) );
  and2f U682 ( .A1(n819), .A2(n818), .Z(n822) );
  or2f U683 ( .A1(n634), .A2(n523), .Z(n542) );
  inv1f U684 ( .I(n1021), .ZN(n1019) );
  and2f U685 ( .A1(n797), .A2(n798), .Z(n582) );
  or2f U686 ( .A1(n795), .A2(n794), .Z(n797) );
  or2f U687 ( .A1(n574), .A2(n685), .Z(n1089) );
  or2f U688 ( .A1(n574), .A2(n1166), .Z(n1083) );
  or2f U689 ( .A1(n924), .A2(n925), .Z(n507) );
  or2f U690 ( .A1(n924), .A2(n925), .Z(n928) );
  and2f U691 ( .A1(n976), .A2(d), .Z(n914) );
  and2f U692 ( .A1(n612), .A2(t), .Z(n701) );
  inv1f U693 ( .I(n1068), .ZN(n1066) );
  or2f U694 ( .A1(n822), .A2(n825), .Z(n629) );
  or2f U695 ( .A1(n574), .A2(n580), .Z(n1095) );
  or2f U696 ( .A1(n613), .A2(n580), .Z(n1179) );
  or2f U701 ( .A1(n1151), .A2(n580), .Z(n1152) );
  or2f U702 ( .A1(n1104), .A2(n580), .Z(n601) );
  inv1f U704 ( .I(n639), .ZN(n599) );
  or2f U706 ( .A1(n859), .A2(n858), .Z(n892) );
  or2f U707 ( .A1(n853), .A2(n852), .Z(n856) );
  inv1f U708 ( .I(n569), .ZN(n726) );
  or2f U710 ( .A1(n537), .A2(n534), .Z(n569) );
  and2f U711 ( .A1(n729), .A2(n730), .Z(n546) );
  inv1 U712 ( .I(n918), .ZN(n920) );
  and2f U713 ( .A1(n570), .A2(a), .Z(n915) );
  or2f U715 ( .A1(n1043), .A2(n1044), .Z(n575) );
  or2f U717 ( .A1(n955), .A2(n956), .Z(n958) );
  or2f U720 ( .A1(n1017), .A2(n1016), .Z(n594) );
  or2f U721 ( .A1(n1017), .A2(n1016), .Z(n1036) );
  or2f U722 ( .A1(n685), .A2(n1166), .Z(n1017) );
  and2f U723 ( .A1(n1026), .A2(i), .Z(n526) );
  or2f U724 ( .A1(n684), .A2(n1117), .Z(n1120) );
  or2f U725 ( .A1(n758), .A2(n628), .Z(n627) );
  or2f U726 ( .A1(n1132), .A2(n554), .Z(n583) );
  or2f U727 ( .A1(n1128), .A2(n1129), .Z(n1132) );
  and2f U728 ( .A1(n590), .A2(p), .Z(n851) );
  or2f U729 ( .A1(n1177), .A2(n615), .Z(n1071) );
  and2f U730 ( .A1(n724), .A2(n723), .Z(n727) );
  or2f U732 ( .A1(n720), .A2(n721), .Z(n724) );
  or2f U733 ( .A1(n1193), .A2(n681), .Z(n829) );
  and2f U734 ( .A1(n1079), .A2(r), .Z(n703) );
  or2f U735 ( .A1(n684), .A2(n1167), .Z(n1170) );
  and2f U736 ( .A1(g), .A2(n653), .Z(n841) );
  or2f U737 ( .A1(n848), .A2(n849), .Z(n671) );
  or2f U739 ( .A1(n518), .A2(n1124), .Z(n647) );
  inv1f U740 ( .I(u), .ZN(n597) );
  or2f U741 ( .A1(n827), .A2(n826), .Z(n523) );
  or2f U748 ( .A1(n1193), .A2(n551), .Z(n564) );
  or2f U756 ( .A1(n1146), .A2(a0), .Z(n1150) );
  or2f U757 ( .A1(n518), .A2(n1145), .Z(n1148) );
  or2f U759 ( .A1(n989), .A2(n988), .Z(n1008) );
  or2f U760 ( .A1(n1043), .A2(n987), .Z(n989) );
  or2f U762 ( .A1(n989), .A2(n988), .Z(n516) );
  and2f U763 ( .A1(f), .A2(n573), .Z(n843) );
  or2f U764 ( .A1(n670), .A2(n539), .Z(n980) );
  or2f U765 ( .A1(n508), .A2(n936), .Z(n1159) );
  and2f U766 ( .A1(s), .A2(n1097), .Z(n700) );
  and2f U767 ( .A1(n566), .A2(n1191), .Z(n603) );
  or2f U768 ( .A1(n589), .A2(n898), .Z(n611) );
  or2f U769 ( .A1(n897), .A2(n901), .Z(n589) );
  or2f U770 ( .A1(n519), .A2(n1111), .Z(n1114) );
  or2f U773 ( .A1(n1195), .A2(n541), .Z(n566) );
  or2f U774 ( .A1(n726), .A2(n525), .Z(n729) );
  and2f U775 ( .A1(n891), .A2(n651), .Z(n860) );
  or2f U776 ( .A1(n652), .A2(n607), .Z(n1063) );
  or2f U778 ( .A1(n1043), .A2(n1044), .Z(n652) );
  or2f U779 ( .A1(n1166), .A2(n639), .Z(n607) );
  and2f U780 ( .A1(n1004), .A2(h), .Z(n842) );
  inv1f U781 ( .I(g), .ZN(n1004) );
  or2f U782 ( .A1(n1159), .A2(n621), .Z(n561) );
  or2f U783 ( .A1(n896), .A2(n568), .Z(n567) );
  and2f U784 ( .A1(n553), .A2(n688), .Z(n893) );
  or2f U785 ( .A1(n644), .A2(n1179), .Z(n1182) );
  and2f U786 ( .A1(b), .A2(n964), .Z(n916) );
  or2f U787 ( .A1(n921), .A2(n922), .Z(n948) );
  or2f U788 ( .A1(n684), .A2(n1173), .Z(n654) );
  and2f U789 ( .A1(u), .A2(n649), .Z(n745) );
  and2f U790 ( .A1(c), .A2(n605), .Z(n913) );
  and2f U795 ( .A1(n553), .A2(n683), .Z(n949) );
  or2f U796 ( .A1(n922), .A2(n921), .Z(n683) );
  or2f U798 ( .A1(n652), .A2(n607), .Z(n513) );
  and2f U799 ( .A1(n781), .A2(n509), .Z(n661) );
  or2f U815 ( .A1(n792), .A2(n666), .Z(n665) );
  or2f U816 ( .A1(n789), .A2(n790), .Z(n792) );
  and2f U817 ( .A1(n792), .A2(n666), .Z(n795) );
  or2f U818 ( .A1(n601), .A2(n1103), .Z(n1124) );
  inv1 U820 ( .I(n716), .ZN(n714) );
  and2f U822 ( .A1(n676), .A2(n602), .Z(n681) );
  and2f U823 ( .A1(n566), .A2(n1191), .Z(n503) );
  or2f U824 ( .A1(n681), .A2(n1193), .Z(n1191) );
  and2f U825 ( .A1(n645), .A2(y), .Z(n712) );
  or2f U826 ( .A1(n931), .A2(n533), .Z(n934) );
  or2f U827 ( .A1(n1083), .A2(n1178), .Z(n1086) );
  and2f U828 ( .A1(n507), .A2(n927), .Z(n533) );
  and2f U829 ( .A1(n717), .A2(n517), .Z(n524) );
  or2f U830 ( .A1(n732), .A2(n546), .Z(n632) );
  or2f U831 ( .A1(n644), .A2(n1077), .Z(n1080) );
  or2f U832 ( .A1(n505), .A2(n1193), .Z(n1077) );
  and2f U835 ( .A1(z), .A2(n1135), .Z(n713) );
  and2f U836 ( .A1(n565), .A2(n891), .Z(n894) );
  inv1f U837 ( .I(n892), .ZN(n891) );
  or2f U838 ( .A1(n646), .A2(n1030), .Z(n1033) );
  inv1f U840 ( .I(n611), .ZN(n902) );
  or2f U841 ( .A1(n1132), .A2(n554), .Z(n1151) );
  or2f U842 ( .A1(n745), .A2(n746), .Z(n749) );
  inv1f U843 ( .I(n993), .ZN(n991) );
  and2f U844 ( .A1(n565), .A2(n947), .Z(n950) );
  or2f U848 ( .A1(n890), .A2(n549), .Z(n565) );
  or2f U860 ( .A1(n646), .A2(n990), .Z(n993) );
  and2f U861 ( .A1(n707), .A2(n706), .Z(n708) );
  or2f U863 ( .A1(n656), .A2(n520), .Z(n554) );
  inv1f U866 ( .I(n705), .ZN(n707) );
  or2f U867 ( .A1(n853), .A2(n852), .Z(n562) );
  and2f U868 ( .A1(n923), .A2(n688), .Z(n861) );
  or2f U869 ( .A1(n670), .A2(n539), .Z(n626) );
  or2f U870 ( .A1(n599), .A2(n987), .Z(n670) );
  or2f U871 ( .A1(n558), .A2(n871), .Z(n639) );
  and2f U872 ( .A1(n869), .A2(n868), .Z(n558) );
  or2f U873 ( .A1(n785), .A2(n661), .Z(n680) );
  or2f U874 ( .A1(n1123), .A2(n685), .Z(n1117) );
  or2f U875 ( .A1(n1123), .A2(n1166), .Z(n1111) );
  and2f U878 ( .A1(n930), .A2(n929), .Z(n931) );
  or2f U879 ( .A1(n1160), .A2(n1178), .Z(n1163) );
  or2f U881 ( .A1(n1073), .A2(n1185), .Z(n1074) );
  and2f U882 ( .A1(n600), .A2(w), .Z(n743) );
  or2f U883 ( .A1(n744), .A2(n743), .Z(n748) );
  and2f U888 ( .A1(n1119), .A2(x), .Z(n744) );
  and2f U898 ( .A1(n824), .A2(n825), .Z(n826) );
  or2f U899 ( .A1(n821), .A2(n571), .Z(n824) );
  and2f U900 ( .A1(n830), .A2(n564), .Z(n604) );
  or2f U904 ( .A1(n635), .A2(n541), .Z(n830) );
  inv1f U905 ( .I(n627), .ZN(n760) );
  or2f U907 ( .A1(n644), .A2(n1152), .Z(n1155) );
  and2f U908 ( .A1(n758), .A2(n628), .Z(n761) );
  and2f U909 ( .A1(n764), .A2(n765), .Z(n766) );
  or2f U910 ( .A1(n713), .A2(n712), .Z(n716) );
  or2f U911 ( .A1(n719), .A2(n718), .Z(n788) );
  and2f U912 ( .A1(n717), .A2(n517), .Z(n718) );
  and2f U913 ( .A1(n1130), .A2(n1102), .Z(n540) );
  or2f U914 ( .A1(n800), .A2(n582), .Z(n1130) );
  or2f U926 ( .A1(n886), .A2(n526), .Z(n527) );
  or2f U927 ( .A1(n500), .A2(n1009), .Z(n1012) );
  inv1f U928 ( .I(n621), .ZN(n1043) );
  or2f U929 ( .A1(n961), .A2(n960), .Z(n621) );
  and2f U930 ( .A1(j), .A2(n1020), .Z(n886) );
  or2f U931 ( .A1(n719), .A2(n524), .Z(n667) );
  and2f U932 ( .A1(n811), .A2(n667), .Z(n789) );
  or2f U933 ( .A1(n1196), .A2(n1045), .Z(n1048) );
  or2f U934 ( .A1(n1064), .A2(n962), .Z(n965) );
  or2f U935 ( .A1(n1064), .A2(n968), .Z(n971) );
  or2f U936 ( .A1(n1196), .A2(n1051), .Z(n1054) );
  inv1f U937 ( .I(j), .ZN(n1026) );
  and2f U938 ( .A1(n1026), .A2(i), .Z(n885) );
  and2f U939 ( .A1(n900), .A2(n901), .Z(n535) );
  or2f U940 ( .A1(n898), .A2(n897), .Z(n900) );
  and2f U941 ( .A1(n502), .A2(n501), .Z(n684) );
  or2f U942 ( .A1(n703), .A2(n702), .Z(n706) );
  and2f U943 ( .A1(q), .A2(n619), .Z(n702) );
  and2f U944 ( .A1(n1189), .A2(n830), .Z(n646) );
  or2f U945 ( .A1(n1193), .A2(n551), .Z(n1189) );
  and2f U946 ( .A1(n676), .A2(n602), .Z(n551) );
  and2f U947 ( .A1(n705), .A2(n704), .Z(n709) );
  or2f U948 ( .A1(n700), .A2(n701), .Z(n705) );
  inv1f U949 ( .I(n706), .ZN(n704) );
  and2f U950 ( .A1(n814), .A2(n680), .Z(n512) );
  or2f U953 ( .A1(n519), .A2(n1133), .Z(n1136) );
  or2f U954 ( .A1(n583), .A2(n515), .Z(n1133) );
  or2f U956 ( .A1(n827), .A2(n522), .Z(n630) );
  and2f U957 ( .A1(n747), .A2(n748), .Z(n752) );
  or2f U958 ( .A1(n843), .A2(n591), .Z(n846) );
  and2f U972 ( .A1(n592), .A2(e), .Z(n591) );
  or2f U973 ( .A1(n871), .A2(n870), .Z(n1177) );
  and2f U974 ( .A1(n868), .A2(n869), .Z(n870) );
  or2f U975 ( .A1(n1044), .A2(n1015), .Z(n1016) );
  inv1f U976 ( .I(n1177), .ZN(n1015) );
  and2f U978 ( .A1(n847), .A2(n846), .Z(n848) );
  or2f U979 ( .A1(n785), .A2(n786), .Z(n813) );
  and2f U980 ( .A1(n781), .A2(n509), .Z(n786) );
  or2f U981 ( .A1(n503), .A2(n974), .Z(n977) );
  or2f U982 ( .A1(n503), .A2(n1002), .Z(n1005) );
  and2f U983 ( .A1(n1181), .A2(e0), .Z(n778) );
  or2f U985 ( .A1(n638), .A2(n766), .Z(n548) );
  or2f U986 ( .A1(n760), .A2(n761), .Z(n1187) );
  or2f U987 ( .A1(n760), .A2(n761), .Z(n764) );
  or2f U996 ( .A1(n709), .A2(n708), .Z(n754) );
  or2f U999 ( .A1(n1159), .A2(n685), .Z(n539) );
  or2f U1000 ( .A1(n961), .A2(n506), .Z(n685) );
  and2f U1001 ( .A1(n588), .A2(n543), .Z(n553) );
  or2f U1002 ( .A1(n527), .A2(n889), .Z(n588) );
  or2f U1003 ( .A1(n887), .A2(n545), .Z(n543) );
  inv1f U1004 ( .I(i), .ZN(n1020) );
  and2f U1005 ( .A1(n958), .A2(n959), .Z(n506) );
  or2f U1006 ( .A1(n799), .A2(n800), .Z(n520) );
  and2f U1007 ( .A1(n797), .A2(n798), .Z(n799) );
  inv1f U1008 ( .I(n618), .ZN(n800) );
  and2f U1009 ( .A1(n784), .A2(n783), .Z(n785) );
  or2f U1010 ( .A1(n596), .A2(n794), .Z(n618) );
  and2f U1011 ( .A1(f0), .A2(n1174), .Z(n659) );
  inv1f U1012 ( .I(n1040), .ZN(n1038) );
  and2f U1013 ( .A1(n857), .A2(n562), .Z(n858) );
  inv1f U1017 ( .I(n855), .ZN(n857) );
  or2f U1018 ( .A1(n603), .A2(n1037), .Z(n1040) );
  and2f U1019 ( .A1(n), .A2(n593), .Z(n853) );
  or2f U1020 ( .A1(n639), .A2(n624), .Z(n988) );
  or2f U1022 ( .A1(n508), .A2(n609), .Z(n624) );
  and2f U1023 ( .A1(n920), .A2(n919), .Z(n921) );
  or2f U1035 ( .A1(n916), .A2(n915), .Z(n919) );
  and2f U1036 ( .A1(n947), .A2(n651), .Z(n925) );
  inv1f U1037 ( .I(n948), .ZN(n947) );
  or2f U1040 ( .A1(n848), .A2(n849), .Z(n651) );
  or2f U1041 ( .A1(n1192), .A2(n1057), .Z(n1060) );
  and2f U1043 ( .A1(n1189), .A2(n566), .Z(n500) );
  or2f U1044 ( .A1(n513), .A2(n1194), .Z(n1057) );
  and2f U1046 ( .A1(n854), .A2(n855), .Z(n859) );
  and2f U1047 ( .A1(n643), .A2(m), .Z(n852) );
  or2f U1049 ( .A1(n902), .A2(n1186), .Z(n1166) );
  and2f U1052 ( .A1(n753), .A2(n667), .Z(n721) );
  and2f U1053 ( .A1(n787), .A2(n680), .Z(n790) );
  or2f U1055 ( .A1(n519), .A2(n1105), .Z(n1108) );
  and2f U1058 ( .A1(n502), .A2(n501), .Z(n519) );
  or2f U1063 ( .A1(n584), .A2(n585), .Z(n1105) );
  inv1f U1064 ( .I(n556), .ZN(n1104) );
  and2f U1069 ( .A1(n1130), .A2(n632), .Z(n556) );
  and2f U1070 ( .A1(n714), .A2(n715), .Z(n719) );
  or2f U1071 ( .A1(n659), .A2(n778), .Z(n782) );
  or2f U1072 ( .A1(n659), .A2(n778), .Z(n509) );
  and2f U1073 ( .A1(n811), .A2(n637), .Z(n816) );
  or2f U1074 ( .A1(n550), .A2(n816), .Z(n677) );
  and2f U1075 ( .A1(n830), .A2(n829), .Z(n1064) );
  or2f U1076 ( .A1(n608), .A2(n508), .Z(n538) );
  or2f U1080 ( .A1(n529), .A2(n530), .Z(n608) );
  and2f U1081 ( .A1(n923), .A2(n683), .Z(n924) );
  inv1f U1083 ( .I(n671), .ZN(n923) );
  or2f U1086 ( .A1(n623), .A2(n622), .Z(n658) );
  and2f U1091 ( .A1(n844), .A2(n845), .Z(n849) );
  or2f U1092 ( .A1(n842), .A2(n841), .Z(n845) );
  or2f U1097 ( .A1(n780), .A2(n779), .Z(n783) );
  or2f U1098 ( .A1(n800), .A2(n799), .Z(n634) );
  or2f U1099 ( .A1(n604), .A2(n996), .Z(n999) );
  or2f U1100 ( .A1(n1197), .A2(n1065), .Z(n1068) );
  or2f U1102 ( .A1(n604), .A2(n1024), .Z(n1027) );
  or2f U1103 ( .A1(n1197), .A2(n1018), .Z(n1021) );
  and2f U1107 ( .A1(n814), .A2(n680), .Z(n815) );
  inv1f U1108 ( .I(n812), .ZN(n814) );
  or2f U1109 ( .A1(n518), .A2(n1139), .Z(n1142) );
  or2f U1114 ( .A1(n1166), .A2(n583), .Z(n1139) );
  or2f U1115 ( .A1(n629), .A2(n821), .Z(n675) );
  and2f U1120 ( .A1(n750), .A2(n572), .Z(n528) );
  or2f U1121 ( .A1(n603), .A2(n981), .Z(n984) );
  or2f U1122 ( .A1(n648), .A2(n626), .Z(n981) );
  or2f U1125 ( .A1(n884), .A2(n883), .Z(n887) );
  and2f U1126 ( .A1(n896), .A2(n568), .Z(n897) );
  or2f U1128 ( .A1(n894), .A2(n893), .Z(n896) );
  or2f U1129 ( .A1(n518), .A2(n1089), .Z(n1092) );
  and2f U1134 ( .A1(n1074), .A2(n1075), .Z(n518) );
  and2f U1135 ( .A1(n953), .A2(n617), .Z(n956) );
  or2f U1139 ( .A1(n950), .A2(n949), .Z(n953) );
  and2f U1140 ( .A1(n917), .A2(n918), .Z(n922) );
  or2f U1146 ( .A1(n914), .A2(n913), .Z(n918) );
  inv1f U1147 ( .I(n919), .ZN(n917) );
  or2f U1151 ( .A1(n575), .A2(n1188), .Z(n1075) );
  or2f U1152 ( .A1(n851), .A2(n850), .Z(n855) );
  and2f U1153 ( .A1(n687), .A2(o), .Z(n850) );
  or2f U1154 ( .A1(n1185), .A2(n1073), .Z(n502) );
  or2f U1155 ( .A1(n987), .A2(n1015), .Z(n1073) );
  or2f U1156 ( .A1(n861), .A2(n860), .Z(n863) );
  and2f U1160 ( .A1(n502), .A2(n501), .Z(n644) );
  or2f U1161 ( .A1(n575), .A2(n1188), .Z(n501) );
  or2f U1162 ( .A1(n756), .A2(n755), .Z(n758) );
  and2f U1166 ( .A1(n753), .A2(n637), .Z(n756) );
  and2f U1167 ( .A1(n814), .A2(n674), .Z(n755) );
  or2f U1168 ( .A1(n635), .A2(n1158), .Z(n613) );
  or2f U1172 ( .A1(n634), .A2(n523), .Z(n1158) );
  or2f U1173 ( .A1(n1128), .A2(n641), .Z(n635) );
  inv1f U1174 ( .I(n650), .ZN(n1128) );
  or2f U1178 ( .A1(n1095), .A2(n1178), .Z(n1098) );
  and2f U1179 ( .A1(n1074), .A2(n1075), .Z(n1178) );
  and2f U1180 ( .A1(n787), .A2(n674), .Z(n720) );
  inv1f U1185 ( .I(n788), .ZN(n787) );
  or2f U1186 ( .A1(n1193), .A2(n499), .Z(n574) );
endmodule

