
module alu4_cl ( n, m, l, k, j, i, h, g, f, e, d, c, b, a, v, u, t, s, r, q, p, 
        o );
  input n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output v, u, t, s, r, q, p, o;
  wire   n1386, n1387, n1, n37, n45, n46, n47, n48, n49, n51, n52, n53, n54,
         n55, n56, n61, n62, n109, n113, n114, n166, n224, n225, n226, n227,
         n234, n249, n264, n275, n276, n277, n283, n366, n367, n368, n389,
         n390, n391, n392, n393, n394, n415, n416, n417, n497, n498, n499,
         n516, n559, n560, n561, n562, n597, n598, n599, n600, n601, n602,
         n662, n663, n701, n702, n703, n704, n705, n706, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395;

  and2 U1 ( .A1(n1), .A2(n1387), .Z(v) );
  and2 U27 ( .A1(n45), .A2(l), .Z(n37) );
  or2 U28 ( .A1(n46), .A2(n47), .Z(n45) );
  or2 U29 ( .A1(n48), .A2(n49), .Z(n47) );
  and2 U30 ( .A1(n1382), .A2(n51), .Z(n49) );
  or2 U31 ( .A1(n1386), .A2(n52), .Z(n51) );
  and2 U32 ( .A1(n53), .A2(n54), .Z(n52) );
  and2 U33 ( .A1(n55), .A2(n56), .Z(n48) );
  or2 U36 ( .A1(n61), .A2(n62), .Z(n46) );
  and2 U71 ( .A1(n113), .A2(n114), .Z(n109) );
  or2 U72 ( .A1(d), .A2(n1383), .Z(n114) );
  or2 U73 ( .A1(h), .A2(n1384), .Z(n113) );
  or2 U166 ( .A1(n225), .A2(n226), .Z(n224) );
  and2 U168 ( .A1(n1381), .A2(d), .Z(n225) );
  and2 U175 ( .A1(l), .A2(n1384), .Z(n234) );
  and2 U186 ( .A1(d), .A2(l), .Z(n249) );
  or2 U203 ( .A1(n1386), .A2(n227), .Z(n1387) );
  inv1 U204 ( .I(n53), .ZN(n227) );
  or2 U205 ( .A1(d), .A2(h), .Z(n53) );
  and2 U206 ( .A1(d), .A2(h), .Z(n1386) );
  or2 U210 ( .A1(n276), .A2(n277), .Z(n264) );
  and2 U214 ( .A1(d), .A2(n1383), .Z(n283) );
  and2 U288 ( .A1(n367), .A2(n368), .Z(n366) );
  and2 U310 ( .A1(n390), .A2(n391), .Z(n389) );
  inv1 U311 ( .I(n392), .ZN(n391) );
  and2 U312 ( .A1(n393), .A2(n275), .Z(n392) );
  and2 U313 ( .A1(n394), .A2(n166), .Z(n390) );
  or2 U336 ( .A1(n416), .A2(n417), .Z(n415) );
  and2 U389 ( .A1(l), .A2(c), .Z(n275) );
  and2 U425 ( .A1(n393), .A2(n498), .Z(n497) );
  or2 U426 ( .A1(l), .A2(n499), .Z(n498) );
  or2 U430 ( .A1(a), .A2(b), .Z(n393) );
  or2 U446 ( .A1(i), .A2(l), .Z(n516) );
  or2 U494 ( .A1(n560), .A2(n561), .Z(n559) );
  and2 U495 ( .A1(n1381), .A2(b), .Z(n561) );
  and2 U496 ( .A1(f), .A2(n562), .Z(n560) );
  or2 U545 ( .A1(n597), .A2(n598), .Z(o) );
  or2 U546 ( .A1(n599), .A2(n600), .Z(n598) );
  or2 U547 ( .A1(n601), .A2(n602), .Z(n600) );
  and2 U602 ( .A1(n1385), .A2(e), .Z(n601) );
  or2 U626 ( .A1(n662), .A2(n663), .Z(n597) );
  and2 U713 ( .A1(n886), .A2(n705), .Z(n704) );
  inv1 U714 ( .I(n888), .ZN(n705) );
  and2 U715 ( .A1(n1180), .A2(n1307), .Z(n706) );
  buf0 U716 ( .I(n1387), .Z(s) );
  buf0 U717 ( .I(n1386), .Z(t) );
  inv1 U720 ( .I(n710), .ZN(n853) );
  or2 U724 ( .A1(n1328), .A2(n1218), .Z(n713) );
  and2 U726 ( .A1(n724), .A2(n717), .Z(n715) );
  or2 U727 ( .A1(n715), .A2(n716), .Z(n718) );
  and2 U728 ( .A1(n1393), .A2(n984), .Z(n716) );
  and2 U729 ( .A1(n1226), .A2(n1393), .Z(n717) );
  inv1 U730 ( .I(n718), .ZN(n720) );
  and2 U735 ( .A1(j), .A2(i), .Z(n722) );
  inv1 U736 ( .I(n722), .ZN(n1368) );
  inv1 U740 ( .I(j), .ZN(n725) );
  inv1 U743 ( .I(i), .ZN(n728) );
  inv1 U744 ( .I(l), .ZN(n729) );
  or2 U745 ( .A1(l), .A2(k), .Z(n761) );
  inv1 U746 ( .I(n), .ZN(n1328) );
  or2 U747 ( .A1(n761), .A2(n1328), .Z(n730) );
  or2 U749 ( .A1(n730), .A2(n1368), .Z(n731) );
  inv1 U750 ( .I(n731), .ZN(n1349) );
  inv1 U751 ( .I(a), .ZN(n1085) );
  or2 U752 ( .A1(n1085), .A2(n745), .Z(n1059) );
  inv1 U753 ( .I(n1059), .ZN(n1062) );
  inv1 U754 ( .I(l), .ZN(n1371) );
  and2 U755 ( .A1(i), .A2(n729), .Z(n732) );
  inv1 U756 ( .I(n761), .ZN(n1308) );
  or2 U757 ( .A1(n732), .A2(n1308), .Z(n734) );
  or2 U758 ( .A1(n), .A2(n725), .Z(n733) );
  or2 U759 ( .A1(n734), .A2(n733), .Z(n735) );
  inv1 U760 ( .I(n735), .ZN(n1342) );
  and2 U761 ( .A1(n1062), .A2(n1342), .Z(n736) );
  or2 U762 ( .A1(n1349), .A2(n736), .Z(n662) );
  inv1 U763 ( .I(k), .ZN(n1205) );
  or2 U764 ( .A1(n940), .A2(n725), .Z(n737) );
  or2 U765 ( .A1(n737), .A2(i), .Z(n833) );
  inv1 U766 ( .I(n833), .ZN(n1029) );
  and2 U767 ( .A1(n1029), .A2(n710), .Z(n748) );
  and2 U768 ( .A1(a), .A2(j), .Z(n738) );
  and2 U769 ( .A1(n738), .A2(n727), .Z(n744) );
  and2 U770 ( .A1(j), .A2(n727), .Z(n739) );
  and2 U771 ( .A1(n940), .A2(n739), .Z(n742) );
  inv1 U773 ( .I(n740), .ZN(n1077) );
  or2 U774 ( .A1(n), .A2(j), .Z(n828) );
  inv1 U775 ( .I(n828), .ZN(n1228) );
  and2 U776 ( .A1(n1077), .A2(n1228), .Z(n741) );
  or2 U777 ( .A1(n742), .A2(n741), .Z(n743) );
  or2 U778 ( .A1(n940), .A2(n1368), .Z(n776) );
  inv1 U779 ( .I(n776), .ZN(n979) );
  or2 U780 ( .A1(n743), .A2(n979), .Z(n868) );
  or2 U781 ( .A1(n744), .A2(n868), .Z(n746) );
  inv1 U782 ( .I(e), .ZN(n745) );
  and2 U783 ( .A1(n746), .A2(n745), .Z(n747) );
  or2 U784 ( .A1(n748), .A2(n747), .Z(n752) );
  and2 U785 ( .A1(l), .A2(n1328), .Z(n749) );
  or2 U786 ( .A1(j), .A2(n1362), .Z(n792) );
  or2 U787 ( .A1(n749), .A2(n792), .Z(n950) );
  inv1 U788 ( .I(n950), .ZN(n887) );
  or2 U789 ( .A1(e), .A2(a), .Z(n750) );
  and2 U790 ( .A1(n887), .A2(n750), .Z(n751) );
  or2 U792 ( .A1(k), .A2(i), .Z(n1046) );
  or2 U793 ( .A1(n1046), .A2(n), .Z(n906) );
  or2 U794 ( .A1(a), .A2(n906), .Z(n753) );
  inv1 U795 ( .I(n753), .ZN(n758) );
  or2 U796 ( .A1(j), .A2(i), .Z(n926) );
  and2 U797 ( .A1(n1368), .A2(n926), .Z(n755) );
  or2 U798 ( .A1(n1328), .A2(k), .Z(n754) );
  or2 U799 ( .A1(n755), .A2(n754), .Z(n756) );
  inv1 U800 ( .I(n756), .ZN(n954) );
  or2 U801 ( .A1(n926), .A2(n940), .Z(n780) );
  inv1 U802 ( .I(n780), .ZN(n974) );
  or2 U803 ( .A1(n954), .A2(n974), .Z(n889) );
  and2 U804 ( .A1(n1062), .A2(n889), .Z(n757) );
  or2 U805 ( .A1(n758), .A2(n757), .Z(n759) );
  or2 U807 ( .A1(n1205), .A2(i), .Z(n763) );
  or2 U808 ( .A1(n761), .A2(n1362), .Z(n762) );
  and2 U809 ( .A1(n763), .A2(n762), .Z(n764) );
  or2 U810 ( .A1(n764), .A2(n828), .Z(n765) );
  inv1 U811 ( .I(n765), .ZN(n1332) );
  and2 U812 ( .A1(n1390), .A2(n1332), .Z(n770) );
  and2 U813 ( .A1(n745), .A2(n1228), .Z(n768) );
  or2 U814 ( .A1(n1085), .A2(n729), .Z(n766) );
  inv1 U815 ( .I(n766), .ZN(n1038) );
  or2 U816 ( .A1(n940), .A2(n1362), .Z(n777) );
  inv1 U817 ( .I(n777), .ZN(n1226) );
  or2 U818 ( .A1(n1038), .A2(n1226), .Z(n767) );
  and2 U819 ( .A1(n768), .A2(n767), .Z(n769) );
  or2 U820 ( .A1(n770), .A2(n769), .Z(n773) );
  or2 U821 ( .A1(n1368), .A2(n1205), .Z(n1206) );
  or2 U822 ( .A1(n1206), .A2(n), .Z(n1111) );
  or2 U823 ( .A1(n1111), .A2(n1032), .Z(n771) );
  inv1 U824 ( .I(n771), .ZN(n772) );
  or2 U825 ( .A1(n773), .A2(n772), .Z(n663) );
  or2 U826 ( .A1(n725), .A2(n729), .Z(n774) );
  or2 U827 ( .A1(n774), .A2(i), .Z(n879) );
  or2 U828 ( .A1(n879), .A2(n), .Z(n775) );
  inv1 U829 ( .I(n775), .ZN(n1385) );
  or2 U831 ( .A1(n777), .A2(j), .Z(n977) );
  or2 U832 ( .A1(n977), .A2(n1059), .Z(n778) );
  or2 U836 ( .A1(n782), .A2(n781), .Z(n783) );
  and2 U838 ( .A1(n979), .A2(n1395), .Z(n791) );
  or2 U839 ( .A1(n1046), .A2(n1085), .Z(n785) );
  or2 U840 ( .A1(n785), .A2(j), .Z(n786) );
  inv1 U841 ( .I(n786), .ZN(n788) );
  or2 U842 ( .A1(n1368), .A2(k), .Z(n787) );
  inv1 U843 ( .I(n787), .ZN(n1049) );
  or2 U844 ( .A1(n1049), .A2(n1029), .Z(n1100) );
  or2 U845 ( .A1(n788), .A2(n1100), .Z(n789) );
  and2 U846 ( .A1(n1390), .A2(n789), .Z(n790) );
  or2 U847 ( .A1(n791), .A2(n790), .Z(n821) );
  or2 U848 ( .A1(n792), .A2(k), .Z(n1210) );
  inv1 U849 ( .I(n1210), .ZN(n1382) );
  and2 U850 ( .A1(a), .A2(n1382), .Z(n793) );
  and2 U851 ( .A1(n745), .A2(n793), .Z(n819) );
  or2 U853 ( .A1(n879), .A2(k), .Z(n794) );
  inv1 U854 ( .I(n794), .ZN(n991) );
  and2 U855 ( .A1(n1062), .A2(n991), .Z(n795) );
  or2 U857 ( .A1(n1071), .A2(n1390), .Z(n797) );
  inv1 U858 ( .I(n797), .ZN(n802) );
  inv1 U861 ( .I(n798), .ZN(n799) );
  or2 U862 ( .A1(n800), .A2(n799), .Z(n801) );
  or2 U863 ( .A1(n802), .A2(n801), .Z(n803) );
  and2 U864 ( .A1(n725), .A2(n803), .Z(n806) );
  inv1 U865 ( .I(n1046), .ZN(n1289) );
  or2 U866 ( .A1(n1099), .A2(a), .Z(n807) );
  and2 U867 ( .A1(n1289), .A2(n807), .Z(n804) );
  or2 U868 ( .A1(n804), .A2(l), .Z(n805) );
  inv1 U870 ( .I(n1206), .ZN(n1310) );
  or2 U871 ( .A1(n807), .A2(n1310), .Z(n811) );
  and2 U872 ( .A1(k), .A2(n1390), .Z(n808) );
  and2 U873 ( .A1(n1368), .A2(n808), .Z(n809) );
  or2 U874 ( .A1(n809), .A2(n1085), .Z(n810) );
  and2 U875 ( .A1(n811), .A2(n810), .Z(n815) );
  or2 U876 ( .A1(n1395), .A2(n1046), .Z(n812) );
  inv1 U877 ( .I(n812), .ZN(n813) );
  or2 U878 ( .A1(n813), .A2(n729), .Z(n814) );
  or2 U879 ( .A1(n815), .A2(n814), .Z(n816) );
  inv1 U883 ( .I(n825), .ZN(n822) );
  and2 U886 ( .A1(n), .A2(n1148), .Z(n827) );
  inv1 U887 ( .I(m), .ZN(n824) );
  or2 U888 ( .A1(n825), .A2(n824), .Z(n826) );
  and2 U889 ( .A1(n827), .A2(n826), .Z(n602) );
  and2 U890 ( .A1(n729), .A2(n1046), .Z(n829) );
  or2 U891 ( .A1(n829), .A2(n828), .Z(n830) );
  inv1 U892 ( .I(n830), .ZN(n1334) );
  and2 U893 ( .A1(n1099), .A2(n1334), .Z(n846) );
  or2 U894 ( .A1(n1046), .A2(n1390), .Z(n831) );
  inv1 U895 ( .I(n831), .ZN(n832) );
  or2 U896 ( .A1(n832), .A2(n745), .Z(n837) );
  or2 U897 ( .A1(a), .A2(n833), .Z(n834) );
  inv1 U898 ( .I(n834), .ZN(n835) );
  or2 U899 ( .A1(n835), .A2(e), .Z(n836) );
  and2 U900 ( .A1(n837), .A2(n836), .Z(n843) );
  or2 U901 ( .A1(n1210), .A2(n729), .Z(n1240) );
  or2 U902 ( .A1(n853), .A2(n1240), .Z(n838) );
  inv1 U903 ( .I(n838), .ZN(n841) );
  inv1 U904 ( .I(n926), .ZN(n1302) );
  or2 U905 ( .A1(n1302), .A2(k), .Z(n1004) );
  inv1 U906 ( .I(n1004), .ZN(n839) );
  or2 U907 ( .A1(n839), .A2(n729), .Z(n876) );
  and2 U908 ( .A1(n1381), .A2(a), .Z(n840) );
  or2 U909 ( .A1(n841), .A2(n840), .Z(n842) );
  or2 U910 ( .A1(n843), .A2(n842), .Z(n844) );
  and2 U911 ( .A1(n844), .A2(n1328), .Z(n845) );
  or2 U912 ( .A1(n846), .A2(n845), .Z(n599) );
  inv1 U914 ( .I(n1240), .ZN(n1142) );
  and2 U915 ( .A1(n1087), .A2(n1142), .Z(n875) );
  or2 U916 ( .A1(b), .A2(n906), .Z(n847) );
  inv1 U917 ( .I(n847), .ZN(n865) );
  and2 U919 ( .A1(n723), .A2(n710), .Z(n849) );
  or2 U921 ( .A1(n1087), .A2(n1025), .Z(n848) );
  inv1 U922 ( .I(n848), .ZN(n1121) );
  and2 U923 ( .A1(n849), .A2(n1121), .Z(n862) );
  and2 U926 ( .A1(n723), .A2(n1063), .Z(n851) );
  or2 U927 ( .A1(n710), .A2(n851), .Z(n852) );
  inv1 U929 ( .I(n891), .ZN(n1064) );
  or2 U931 ( .A1(b), .A2(f), .Z(n1057) );
  inv1 U932 ( .I(n1057), .ZN(n1028) );
  or2 U933 ( .A1(n853), .A2(n1028), .Z(n854) );
  or2 U936 ( .A1(n729), .A2(n1205), .Z(n857) );
  inv1 U937 ( .I(n857), .ZN(n928) );
  and2 U938 ( .A1(a), .A2(n928), .Z(n858) );
  or2 U939 ( .A1(j), .A2(n858), .Z(n859) );
  or2 U941 ( .A1(n862), .A2(n861), .Z(n863) );
  and2 U942 ( .A1(n727), .A2(n863), .Z(n864) );
  or2 U943 ( .A1(n865), .A2(n864), .Z(n867) );
  and2 U944 ( .A1(n889), .A2(n1121), .Z(n866) );
  and2 U946 ( .A1(n887), .A2(n1057), .Z(n871) );
  inv1 U947 ( .I(n868), .ZN(n949) );
  or2 U948 ( .A1(f), .A2(n949), .Z(n869) );
  inv1 U949 ( .I(n869), .ZN(n870) );
  or2 U950 ( .A1(n871), .A2(n870), .Z(n872) );
  and2 U952 ( .A1(n1289), .A2(n1393), .Z(n874) );
  or2 U953 ( .A1(n875), .A2(n874), .Z(n562) );
  inv1 U954 ( .I(n876), .ZN(n1381) );
  and2 U955 ( .A1(b), .A2(j), .Z(n877) );
  or2 U956 ( .A1(n877), .A2(n1121), .Z(n878) );
  and2 U957 ( .A1(n1226), .A2(n878), .Z(n880) );
  inv1 U958 ( .I(n879), .ZN(n973) );
  or2 U959 ( .A1(n880), .A2(n973), .Z(n881) );
  and2 U960 ( .A1(n1392), .A2(n881), .Z(n883) );
  and2 U963 ( .A1(n1395), .A2(n721), .Z(n885) );
  inv1 U964 ( .I(n1395), .ZN(n921) );
  and2 U965 ( .A1(n921), .A2(n724), .Z(n884) );
  or2 U966 ( .A1(n885), .A2(n884), .Z(n499) );
  or2 U967 ( .A1(c), .A2(g), .Z(n1006) );
  inv1 U968 ( .I(n1006), .ZN(n1016) );
  and2 U969 ( .A1(n1029), .A2(n1016), .Z(n416) );
  and2 U970 ( .A1(n275), .A2(n1004), .Z(n417) );
  or2 U971 ( .A1(n949), .A2(g), .Z(n886) );
  and2 U972 ( .A1(n887), .A2(n1006), .Z(n888) );
  inv1 U973 ( .I(c), .ZN(n1180) );
  inv1 U974 ( .I(g), .ZN(n1131) );
  or2 U975 ( .A1(n1180), .A2(n1131), .Z(n935) );
  inv1 U976 ( .I(n935), .ZN(n1140) );
  and2 U977 ( .A1(n889), .A2(n1140), .Z(n911) );
  and2 U978 ( .A1(b), .A2(n928), .Z(n890) );
  or2 U979 ( .A1(n890), .A2(j), .Z(n901) );
  or2 U980 ( .A1(n1180), .A2(g), .Z(n961) );
  inv1 U981 ( .I(n961), .ZN(n895) );
  or2 U982 ( .A1(c), .A2(n1131), .Z(n932) );
  inv1 U983 ( .I(n932), .ZN(n1141) );
  or2 U988 ( .A1(n895), .A2(n894), .Z(n898) );
  inv1 U989 ( .I(n959), .ZN(n896) );
  or2 U990 ( .A1(n896), .A2(n1016), .Z(n897) );
  and2 U991 ( .A1(n898), .A2(n897), .Z(n899) );
  or2 U992 ( .A1(n899), .A2(n725), .Z(n900) );
  and2 U994 ( .A1(n723), .A2(n1140), .Z(n902) );
  and2 U995 ( .A1(n902), .A2(n959), .Z(n903) );
  or2 U996 ( .A1(n904), .A2(n903), .Z(n905) );
  and2 U997 ( .A1(n727), .A2(n905), .Z(n909) );
  or2 U998 ( .A1(n906), .A2(c), .Z(n907) );
  inv1 U999 ( .I(n907), .ZN(n908) );
  or2 U1000 ( .A1(n909), .A2(n908), .Z(n910) );
  or2 U1001 ( .A1(n911), .A2(n910), .Z(n912) );
  and2 U1003 ( .A1(c), .A2(j), .Z(n913) );
  or2 U1004 ( .A1(n913), .A2(n1140), .Z(n914) );
  and2 U1005 ( .A1(n1226), .A2(n914), .Z(n916) );
  or2 U1007 ( .A1(n916), .A2(n915), .Z(n917) );
  and2 U1009 ( .A1(c), .A2(n973), .Z(n919) );
  or2 U1012 ( .A1(n922), .A2(n721), .Z(n1246) );
  and2 U1014 ( .A1(n1395), .A2(n724), .Z(n923) );
  or2 U1015 ( .A1(n1196), .A2(n923), .Z(n924) );
  or2 U1018 ( .A1(c), .A2(n393), .Z(n166) );
  or2 U1019 ( .A1(n926), .A2(n729), .Z(n927) );
  inv1 U1020 ( .I(n927), .ZN(n930) );
  and2 U1021 ( .A1(n1368), .A2(n928), .Z(n929) );
  or2 U1022 ( .A1(n930), .A2(n929), .Z(n1307) );
  and2 U1023 ( .A1(n1062), .A2(n1057), .Z(n931) );
  or2 U1024 ( .A1(n931), .A2(n1121), .Z(n1005) );
  and2 U1025 ( .A1(n932), .A2(n961), .Z(n933) );
  or2 U1026 ( .A1(n1005), .A2(n933), .Z(n367) );
  or2 U1027 ( .A1(n1006), .A2(n729), .Z(n934) );
  and2 U1028 ( .A1(n935), .A2(n934), .Z(n937) );
  inv1 U1029 ( .I(n1005), .ZN(n936) );
  or2 U1030 ( .A1(n937), .A2(n936), .Z(n368) );
  inv1 U1031 ( .I(h), .ZN(n1383) );
  or2 U1032 ( .A1(n), .A2(d), .Z(n938) );
  or2 U1033 ( .A1(n938), .A2(k), .Z(n939) );
  inv1 U1034 ( .I(n939), .ZN(n276) );
  and2 U1035 ( .A1(n959), .A2(n961), .Z(n945) );
  inv1 U1036 ( .I(n283), .ZN(n943) );
  or2 U1037 ( .A1(n1383), .A2(d), .Z(n941) );
  or2 U1038 ( .A1(n941), .A2(n940), .Z(n942) );
  and2 U1039 ( .A1(n943), .A2(n942), .Z(n944) );
  or2 U1040 ( .A1(n945), .A2(n944), .Z(n947) );
  or2 U1041 ( .A1(n1141), .A2(n725), .Z(n946) );
  or2 U1042 ( .A1(n947), .A2(n946), .Z(n948) );
  inv1 U1043 ( .I(n948), .ZN(n277) );
  inv1 U1044 ( .I(d), .ZN(n1384) );
  and2 U1045 ( .A1(n227), .A2(n1029), .Z(n226) );
  or2 U1046 ( .A1(n949), .A2(h), .Z(n952) );
  or2 U1047 ( .A1(n950), .A2(n227), .Z(n951) );
  and2 U1048 ( .A1(n952), .A2(n951), .Z(n953) );
  inv1 U1049 ( .I(n953), .ZN(n972) );
  and2 U1050 ( .A1(n725), .A2(n723), .Z(n955) );
  or2 U1051 ( .A1(n955), .A2(n954), .Z(n956) );
  and2 U1052 ( .A1(n1386), .A2(n956), .Z(n970) );
  and2 U1053 ( .A1(n1387), .A2(j), .Z(n957) );
  and2 U1054 ( .A1(n723), .A2(n957), .Z(n963) );
  or2 U1055 ( .A1(n1141), .A2(n959), .Z(n960) );
  and2 U1056 ( .A1(n961), .A2(n960), .Z(n962) );
  and2 U1057 ( .A1(n963), .A2(n962), .Z(n964) );
  or2 U1058 ( .A1(n964), .A2(n264), .Z(n965) );
  and2 U1060 ( .A1(n275), .A2(k), .Z(n966) );
  and2 U1061 ( .A1(n1302), .A2(n966), .Z(n967) );
  or2 U1062 ( .A1(n968), .A2(n967), .Z(n969) );
  or2 U1065 ( .A1(n1333), .A2(d), .Z(n56) );
  and2 U1066 ( .A1(n56), .A2(n973), .Z(n976) );
  and2 U1068 ( .A1(n974), .A2(n1335), .Z(n975) );
  or2 U1069 ( .A1(n976), .A2(n975), .Z(n983) );
  inv1 U1070 ( .I(n977), .ZN(n1272) );
  and2 U1071 ( .A1(n1386), .A2(n1272), .Z(n981) );
  or2 U1072 ( .A1(n1335), .A2(n1384), .Z(n978) );
  inv1 U1073 ( .I(n978), .ZN(n1347) );
  and2 U1074 ( .A1(n979), .A2(n1347), .Z(n980) );
  and2 U1077 ( .A1(n1226), .A2(n724), .Z(n985) );
  and2 U1078 ( .A1(n991), .A2(n1121), .Z(n984) );
  inv1 U1080 ( .I(n1197), .ZN(n1079) );
  and2 U1082 ( .A1(n991), .A2(n1140), .Z(n986) );
  and2 U1083 ( .A1(n1079), .A2(n709), .Z(n989) );
  and2 U1084 ( .A1(n1071), .A2(n721), .Z(n1198) );
  inv1 U1085 ( .I(n1198), .ZN(n988) );
  and2 U1086 ( .A1(n989), .A2(n988), .Z(n990) );
  or2 U1087 ( .A1(n990), .A2(n1196), .Z(n1291) );
  inv1 U1088 ( .I(n1291), .ZN(n1287) );
  and2 U1091 ( .A1(n1386), .A2(n991), .Z(n992) );
  or2 U1093 ( .A1(n1287), .A2(n1284), .Z(n994) );
  and2 U1094 ( .A1(n1358), .A2(n994), .Z(n61) );
  or2 U1095 ( .A1(n166), .A2(d), .Z(n995) );
  or2 U1096 ( .A1(n995), .A2(n1206), .Z(n996) );
  inv1 U1097 ( .I(n996), .ZN(n62) );
  and2 U1098 ( .A1(n1180), .A2(n701), .Z(n1002) );
  and2 U1099 ( .A1(n1087), .A2(n1032), .Z(n999) );
  or2 U1100 ( .A1(n1032), .A2(n1087), .Z(n997) );
  and2 U1101 ( .A1(n1391), .A2(n997), .Z(n998) );
  or2 U1102 ( .A1(n999), .A2(n998), .Z(n1159) );
  or2 U1103 ( .A1(n701), .A2(n1180), .Z(n1000) );
  and2 U1104 ( .A1(n1159), .A2(n1000), .Z(n1001) );
  or2 U1105 ( .A1(n1002), .A2(n1001), .Z(n1297) );
  inv1 U1106 ( .I(n1297), .ZN(n1296) );
  or2 U1107 ( .A1(n1296), .A2(n1347), .Z(n1003) );
  and2 U1108 ( .A1(n1004), .A2(n1003), .Z(n55) );
  and2 U1109 ( .A1(n1006), .A2(n1005), .Z(n1007) );
  or2 U1110 ( .A1(n1007), .A2(n1140), .Z(n54) );
  and2 U1111 ( .A1(n1121), .A2(n1016), .Z(n1009) );
  or2 U1112 ( .A1(n1028), .A2(n1121), .Z(n1018) );
  and2 U1113 ( .A1(n1140), .A2(n1018), .Z(n1008) );
  or2 U1114 ( .A1(n1009), .A2(n1008), .Z(n1010) );
  and2 U1115 ( .A1(n1085), .A2(n1010), .Z(n1014) );
  or2 U1116 ( .A1(n166), .A2(f), .Z(n1011) );
  or2 U1117 ( .A1(n1011), .A2(g), .Z(n1012) );
  inv1 U1118 ( .I(n1012), .ZN(n1013) );
  or2 U1119 ( .A1(n1014), .A2(n1013), .Z(n1015) );
  and2 U1120 ( .A1(n745), .A2(n1015), .Z(n1021) );
  or2 U1121 ( .A1(n1140), .A2(n1016), .Z(n1017) );
  and2 U1122 ( .A1(n1062), .A2(n1017), .Z(n1019) );
  and2 U1123 ( .A1(n1019), .A2(n1018), .Z(n1020) );
  or2 U1124 ( .A1(n1021), .A2(n1020), .Z(n1) );
  and2 U1125 ( .A1(b), .A2(l), .Z(n1022) );
  or2 U1126 ( .A1(n1022), .A2(n1226), .Z(n1023) );
  and2 U1127 ( .A1(n1228), .A2(n1023), .Z(n1024) );
  or2 U1128 ( .A1(n1024), .A2(f), .Z(n1027) );
  or2 U1129 ( .A1(n1385), .A2(n1025), .Z(n1026) );
  and2 U1130 ( .A1(n1027), .A2(n1026), .Z(n1120) );
  and2 U1131 ( .A1(n1029), .A2(n1028), .Z(n1030) );
  or2 U1132 ( .A1(n1030), .A2(n559), .Z(n1031) );
  or2 U1133 ( .A1(n1031), .A2(n), .Z(n1110) );
  and2 U1134 ( .A1(n719), .A2(n1393), .Z(n1034) );
  and2 U1135 ( .A1(n1032), .A2(n1391), .Z(n1033) );
  or2 U1136 ( .A1(n1034), .A2(n1033), .Z(n1037) );
  inv1 U1137 ( .I(n1037), .ZN(n1035) );
  and2 U1138 ( .A1(n1307), .A2(n1035), .Z(n1036) );
  or2 U1139 ( .A1(n1036), .A2(b), .Z(n1044) );
  and2 U1140 ( .A1(n1307), .A2(n1037), .Z(n1040) );
  and2 U1141 ( .A1(n1310), .A2(n1038), .Z(n1039) );
  or2 U1142 ( .A1(n1040), .A2(n1039), .Z(n1042) );
  or2 U1143 ( .A1(n1308), .A2(n1087), .Z(n1041) );
  or2 U1144 ( .A1(n1042), .A2(n1041), .Z(n1043) );
  and2 U1145 ( .A1(n1044), .A2(n1043), .Z(n1056) );
  inv1 U1146 ( .I(n497), .ZN(n1045) );
  and2 U1147 ( .A1(n1045), .A2(n1310), .Z(n1054) );
  or2 U1148 ( .A1(n1046), .A2(l), .Z(n1047) );
  inv1 U1149 ( .I(n1047), .ZN(n1052) );
  inv1 U1150 ( .I(n516), .ZN(n1048) );
  and2 U1151 ( .A1(n1048), .A2(j), .Z(n1050) );
  or2 U1152 ( .A1(n1050), .A2(n1049), .Z(n1275) );
  and2 U1153 ( .A1(n1099), .A2(n1275), .Z(n1051) );
  or2 U1154 ( .A1(n1052), .A2(n1051), .Z(n1276) );
  and2 U1155 ( .A1(n1393), .A2(n1276), .Z(n1053) );
  or2 U1156 ( .A1(n1054), .A2(n1053), .Z(n1055) );
  or2 U1157 ( .A1(n1056), .A2(n1055), .Z(n1107) );
  and2 U1158 ( .A1(f), .A2(n729), .Z(n1069) );
  or2 U1159 ( .A1(n1057), .A2(n729), .Z(n1058) );
  inv1 U1160 ( .I(n1058), .ZN(n1061) );
  or2 U1161 ( .A1(n1121), .A2(n1059), .Z(n1060) );
  or2 U1162 ( .A1(n1061), .A2(n1060), .Z(n1067) );
  or2 U1163 ( .A1(n1063), .A2(n1062), .Z(n1065) );
  or2 U1164 ( .A1(n1065), .A2(n1064), .Z(n1066) );
  and2 U1165 ( .A1(n1067), .A2(n1066), .Z(n1068) );
  or2 U1166 ( .A1(n1069), .A2(n1068), .Z(n1070) );
  and2 U1167 ( .A1(n1382), .A2(n1070), .Z(n1076) );
  and2 U1169 ( .A1(n1078), .A2(n721), .Z(n1073) );
  and2 U1170 ( .A1(n1071), .A2(n724), .Z(n1072) );
  or2 U1171 ( .A1(n1073), .A2(n1072), .Z(n1074) );
  and2 U1172 ( .A1(n1205), .A2(n1074), .Z(n1075) );
  or2 U1173 ( .A1(n1076), .A2(n1075), .Z(n1105) );
  and2 U1174 ( .A1(n725), .A2(n1077), .Z(n1084) );
  inv1 U1176 ( .I(n1080), .ZN(n1168) );
  or2 U1177 ( .A1(n1168), .A2(n720), .Z(n1082) );
  or2 U1178 ( .A1(n718), .A2(n1080), .Z(n1081) );
  and2 U1180 ( .A1(n1084), .A2(n1083), .Z(n1097) );
  and2 U1183 ( .A1(b), .A2(n724), .Z(n1089) );
  and2 U1184 ( .A1(n1087), .A2(n721), .Z(n1088) );
  or2 U1185 ( .A1(n1089), .A2(n1088), .Z(n1091) );
  or2 U1186 ( .A1(n1178), .A2(n1091), .Z(n1090) );
  and2 U1187 ( .A1(n1302), .A2(n1090), .Z(n1095) );
  inv1 U1188 ( .I(n1091), .ZN(n1092) );
  or2 U1189 ( .A1(n1093), .A2(n1092), .Z(n1094) );
  and2 U1190 ( .A1(n1095), .A2(n1094), .Z(n1096) );
  or2 U1193 ( .A1(n1393), .A2(n1099), .Z(n1102) );
  inv1 U1194 ( .I(n1100), .ZN(n1101) );
  or2 U1195 ( .A1(n1102), .A2(n1101), .Z(n1318) );
  inv1 U1196 ( .I(n1318), .ZN(n1154) );
  or2 U1197 ( .A1(n1103), .A2(n1154), .Z(n1104) );
  or2 U1201 ( .A1(n1108), .A2(n1328), .Z(n1109) );
  and2 U1202 ( .A1(n1110), .A2(n1109), .Z(n1118) );
  or2 U1203 ( .A1(n1393), .A2(n1332), .Z(n1116) );
  inv1 U1204 ( .I(n1111), .ZN(n1348) );
  and2 U1205 ( .A1(b), .A2(n1348), .Z(n1114) );
  or2 U1206 ( .A1(n1391), .A2(n1334), .Z(n1113) );
  or2 U1207 ( .A1(n1114), .A2(n1113), .Z(n1115) );
  and2 U1208 ( .A1(n1116), .A2(n1115), .Z(n1117) );
  or2 U1209 ( .A1(n1118), .A2(n1117), .Z(n1119) );
  or2 U1210 ( .A1(n1120), .A2(n1119), .Z(n1128) );
  and2 U1211 ( .A1(n1342), .A2(n1121), .Z(n1126) );
  inv1 U1212 ( .I(n1148), .ZN(n1123) );
  and2 U1214 ( .A1(n1123), .A2(n1149), .Z(n1124) );
  or2 U1215 ( .A1(n1124), .A2(n1349), .Z(n1125) );
  or2 U1216 ( .A1(n1126), .A2(n1125), .Z(n1127) );
  or2 U1217 ( .A1(n1128), .A2(n1127), .Z(p) );
  or2 U1218 ( .A1(n1226), .A2(n275), .Z(n1129) );
  and2 U1219 ( .A1(n1228), .A2(n1129), .Z(n1130) );
  or2 U1220 ( .A1(n1130), .A2(g), .Z(n1133) );
  or2 U1221 ( .A1(n1385), .A2(n1131), .Z(n1132) );
  and2 U1222 ( .A1(n1133), .A2(n1132), .Z(n1139) );
  or2 U1223 ( .A1(n1317), .A2(n1332), .Z(n1137) );
  and2 U1224 ( .A1(c), .A2(n1348), .Z(n1135) );
  or2 U1225 ( .A1(n701), .A2(n1334), .Z(n1134) );
  or2 U1226 ( .A1(n1135), .A2(n1134), .Z(n1136) );
  and2 U1227 ( .A1(n1137), .A2(n1136), .Z(n1138) );
  or2 U1228 ( .A1(n1139), .A2(n1138), .Z(n1225) );
  and2 U1229 ( .A1(n1342), .A2(n1140), .Z(n1223) );
  and2 U1230 ( .A1(n1142), .A2(n1141), .Z(n1143) );
  or2 U1231 ( .A1(n1143), .A2(n415), .Z(n1147) );
  and2 U1232 ( .A1(g), .A2(n1289), .Z(n1144) );
  and2 U1233 ( .A1(n1317), .A2(n1144), .Z(n1145) );
  or2 U1234 ( .A1(n1145), .A2(n), .Z(n1146) );
  or2 U1235 ( .A1(n1147), .A2(n1146), .Z(n1220) );
  inv1 U1237 ( .I(n1327), .ZN(n1216) );
  or2 U1238 ( .A1(n701), .A2(n1276), .Z(n1153) );
  and2 U1239 ( .A1(n1393), .A2(n1275), .Z(n1151) );
  and2 U1240 ( .A1(n706), .A2(n1159), .Z(n1150) );
  or2 U1241 ( .A1(n1151), .A2(n1150), .Z(n1152) );
  or2 U1242 ( .A1(n1153), .A2(n1152), .Z(n1158) );
  or2 U1243 ( .A1(n1317), .A2(n1154), .Z(n1156) );
  inv1 U1244 ( .I(n1159), .ZN(n1160) );
  and2 U1245 ( .A1(n706), .A2(n1160), .Z(n1155) );
  or2 U1246 ( .A1(n1156), .A2(n1155), .Z(n1157) );
  and2 U1247 ( .A1(n1158), .A2(n1157), .Z(n1167) );
  and2 U1248 ( .A1(n701), .A2(n1159), .Z(n1162) );
  and2 U1249 ( .A1(n1317), .A2(n1160), .Z(n1161) );
  or2 U1250 ( .A1(n1162), .A2(n1161), .Z(n1163) );
  and2 U1251 ( .A1(n1307), .A2(n1163), .Z(n1164) );
  or2 U1252 ( .A1(n1308), .A2(n1164), .Z(n1165) );
  and2 U1253 ( .A1(c), .A2(n1165), .Z(n1166) );
  or2 U1254 ( .A1(n1167), .A2(n1166), .Z(n1195) );
  inv1 U1257 ( .I(n1265), .ZN(n1170) );
  inv1 U1261 ( .I(n1174), .ZN(n1173) );
  and2 U1262 ( .A1(n703), .A2(n1173), .Z(n1176) );
  and2 U1263 ( .A1(n709), .A2(n1174), .Z(n1175) );
  and2 U1266 ( .A1(b), .A2(n721), .Z(n1179) );
  or2 U1270 ( .A1(n1182), .A2(n1181), .Z(n1185) );
  and2 U1272 ( .A1(n1250), .A2(n1183), .Z(n1187) );
  inv1 U1273 ( .I(n1250), .ZN(n1184) );
  and2 U1274 ( .A1(n1185), .A2(n1184), .Z(n1186) );
  or2 U1275 ( .A1(n1187), .A2(n1186), .Z(n1188) );
  and2 U1276 ( .A1(n1302), .A2(n1188), .Z(n1190) );
  and2 U1277 ( .A1(g), .A2(n1382), .Z(n1189) );
  or2 U1278 ( .A1(n1190), .A2(n1189), .Z(n1191) );
  or2 U1283 ( .A1(n1198), .A2(n1197), .Z(n1199) );
  and2 U1284 ( .A1(n1200), .A2(n1199), .Z(n1203) );
  or2 U1285 ( .A1(n1200), .A2(n1199), .Z(n1201) );
  inv1 U1286 ( .I(n1201), .ZN(n1202) );
  or2 U1287 ( .A1(n1203), .A2(n1202), .Z(n1204) );
  and2 U1288 ( .A1(n1205), .A2(n1204), .Z(n1209) );
  or2 U1289 ( .A1(n389), .A2(n1206), .Z(n1207) );
  inv1 U1290 ( .I(n1207), .ZN(n1208) );
  or2 U1291 ( .A1(n1209), .A2(n1208), .Z(n1213) );
  or2 U1292 ( .A1(n366), .A2(n1210), .Z(n1211) );
  inv1 U1293 ( .I(n1211), .ZN(n1212) );
  or2 U1302 ( .A1(n1226), .A2(n249), .Z(n1227) );
  and2 U1303 ( .A1(n1228), .A2(n1227), .Z(n1229) );
  or2 U1304 ( .A1(n1229), .A2(h), .Z(n1231) );
  or2 U1305 ( .A1(n1385), .A2(n1383), .Z(n1230) );
  and2 U1306 ( .A1(n1231), .A2(n1230), .Z(n1341) );
  and2 U1307 ( .A1(n234), .A2(n1382), .Z(n1233) );
  and2 U1308 ( .A1(n1289), .A2(n1333), .Z(n1232) );
  or2 U1309 ( .A1(n1233), .A2(n1232), .Z(n1234) );
  and2 U1310 ( .A1(h), .A2(n1234), .Z(n1235) );
  or2 U1311 ( .A1(n1235), .A2(n224), .Z(n1236) );
  or2 U1312 ( .A1(n1236), .A2(n), .Z(n1331) );
  inv1 U1313 ( .I(n109), .ZN(n1237) );
  and2 U1314 ( .A1(n1237), .A2(n1382), .Z(n1238) );
  or2 U1315 ( .A1(n1238), .A2(n54), .Z(n1244) );
  inv1 U1316 ( .I(n1387), .ZN(n1239) );
  or2 U1317 ( .A1(n1240), .A2(n1239), .Z(n1241) );
  and2 U1318 ( .A1(n54), .A2(n1241), .Z(n1242) );
  inv1 U1319 ( .I(n1242), .ZN(n1243) );
  and2 U1320 ( .A1(n1244), .A2(n1243), .Z(n1263) );
  and2 U1321 ( .A1(h), .A2(n1382), .Z(n1260) );
  and2 U1323 ( .A1(n1310), .A2(n1245), .Z(n1248) );
  inv1 U1324 ( .I(n1246), .ZN(n1369) );
  or2 U1325 ( .A1(n1358), .A2(n1369), .Z(n1247) );
  and2 U1326 ( .A1(n1248), .A2(n1247), .Z(n1258) );
  and2 U1331 ( .A1(n1370), .A2(n1359), .Z(n1253) );
  or2 U1332 ( .A1(n1254), .A2(n1253), .Z(n1301) );
  inv1 U1333 ( .I(n1301), .ZN(n1256) );
  and2 U1334 ( .A1(d), .A2(n1302), .Z(n1255) );
  and2 U1335 ( .A1(n1256), .A2(n1255), .Z(n1257) );
  or2 U1336 ( .A1(n1258), .A2(n1257), .Z(n1259) );
  or2 U1341 ( .A1(n1266), .A2(n1265), .Z(n1363) );
  inv1 U1342 ( .I(n1284), .ZN(n1283) );
  or2 U1343 ( .A1(n1283), .A2(n1335), .Z(n1267) );
  inv1 U1344 ( .I(n1267), .ZN(n1365) );
  and2 U1345 ( .A1(n1363), .A2(n1365), .Z(n1270) );
  inv1 U1346 ( .I(n1363), .ZN(n1268) );
  and2 U1347 ( .A1(n1268), .A2(n1267), .Z(n1269) );
  or2 U1348 ( .A1(n1270), .A2(n1269), .Z(n1271) );
  and2 U1349 ( .A1(n1272), .A2(n1271), .Z(n1280) );
  or2 U1350 ( .A1(n1317), .A2(n1393), .Z(n1274) );
  and2 U1351 ( .A1(n1275), .A2(n1274), .Z(n1277) );
  or2 U1352 ( .A1(n1277), .A2(n1276), .Z(n1278) );
  and2 U1353 ( .A1(n1333), .A2(n1278), .Z(n1279) );
  or2 U1354 ( .A1(n1280), .A2(n1279), .Z(n1281) );
  and2 U1356 ( .A1(n1358), .A2(n1283), .Z(n1286) );
  and2 U1357 ( .A1(n1370), .A2(n1284), .Z(n1285) );
  or2 U1358 ( .A1(n1286), .A2(n1285), .Z(n1290) );
  or2 U1359 ( .A1(n1290), .A2(n1287), .Z(n1288) );
  inv1 U1361 ( .I(n1290), .ZN(n1292) );
  or2 U1362 ( .A1(n1292), .A2(n1291), .Z(n1293) );
  and2 U1363 ( .A1(n1294), .A2(n1293), .Z(n1295) );
  and2 U1365 ( .A1(n1333), .A2(n1296), .Z(n1299) );
  and2 U1366 ( .A1(n1335), .A2(n1297), .Z(n1298) );
  or2 U1367 ( .A1(n1299), .A2(n1298), .Z(n1306) );
  inv1 U1368 ( .I(n1306), .ZN(n1300) );
  and2 U1369 ( .A1(n1307), .A2(n1300), .Z(n1305) );
  and2 U1370 ( .A1(n1302), .A2(n1301), .Z(n1303) );
  or2 U1371 ( .A1(n1303), .A2(d), .Z(n1304) );
  or2 U1372 ( .A1(n1305), .A2(n1304), .Z(n1316) );
  and2 U1373 ( .A1(n1307), .A2(n1306), .Z(n1309) );
  or2 U1374 ( .A1(n1309), .A2(n1308), .Z(n1314) );
  and2 U1375 ( .A1(l), .A2(n1310), .Z(n1311) );
  and2 U1376 ( .A1(n166), .A2(n1311), .Z(n1312) );
  or2 U1377 ( .A1(n1312), .A2(n1384), .Z(n1313) );
  or2 U1378 ( .A1(n1314), .A2(n1313), .Z(n1315) );
  and2 U1379 ( .A1(n1316), .A2(n1315), .Z(n1321) );
  or2 U1380 ( .A1(n1318), .A2(n1317), .Z(n1319) );
  or2 U1381 ( .A1(n1319), .A2(n1333), .Z(n1320) );
  inv1 U1382 ( .I(n1320), .ZN(n1374) );
  or2 U1383 ( .A1(n1321), .A2(n1374), .Z(n1322) );
  or2 U1390 ( .A1(n1333), .A2(n1332), .Z(n1337) );
  or2 U1391 ( .A1(n1335), .A2(n1334), .Z(n1336) );
  and2 U1392 ( .A1(n1337), .A2(n1336), .Z(n1338) );
  and2 U1395 ( .A1(n1386), .A2(n1342), .Z(n1346) );
  inv1 U1396 ( .I(n1356), .ZN(n1344) );
  inv1 U1397 ( .I(n1343), .ZN(n1355) );
  and2 U1398 ( .A1(n1344), .A2(n1355), .Z(n1345) );
  or2 U1399 ( .A1(n1346), .A2(n1345), .Z(n1352) );
  and2 U1400 ( .A1(n1348), .A2(n1347), .Z(n1350) );
  or2 U1401 ( .A1(n1350), .A2(n1349), .Z(n1351) );
  or2 U1402 ( .A1(n1352), .A2(n1351), .Z(n1353) );
  or2 U1403 ( .A1(n1354), .A2(n1353), .Z(r) );
  or2 U1405 ( .A1(n1357), .A2(n37), .Z(n1379) );
  and2 U1406 ( .A1(d), .A2(n1358), .Z(n1360) );
  or2 U1407 ( .A1(n1360), .A2(n1359), .Z(n1361) );
  and2 U1408 ( .A1(n1362), .A2(n1361), .Z(n1364) );
  or2 U1409 ( .A1(n1364), .A2(n1363), .Z(n1366) );
  or2 U1410 ( .A1(n1366), .A2(n1365), .Z(n1367) );
  and2 U1411 ( .A1(n725), .A2(n1367), .Z(n1377) );
  and2 U1412 ( .A1(n722), .A2(n1369), .Z(n1373) );
  and2 U1413 ( .A1(n729), .A2(n1370), .Z(n1372) );
  and2 U1414 ( .A1(n1373), .A2(n1372), .Z(n1375) );
  or2 U1415 ( .A1(n1375), .A2(n1374), .Z(n1376) );
  or2 U1416 ( .A1(n1377), .A2(n1376), .Z(n1378) );
  or2 U1417 ( .A1(n1379), .A2(n1378), .Z(n1380) );
  and2 U1418 ( .A1(n), .A2(n1380), .Z(u) );
  or2f U709 ( .A1(n985), .A2(n984), .Z(n1197) );
  inv1f U710 ( .I(n719), .ZN(n1032) );
  and2 U711 ( .A1(n1099), .A2(n879), .Z(n782) );
  or2f U712 ( .A1(n1395), .A2(n1085), .Z(n1093) );
  or2f U718 ( .A1(n1395), .A2(a), .Z(n798) );
  inv1f U719 ( .I(n1394), .ZN(n1395) );
  or2f U721 ( .A1(n796), .A2(n795), .Z(n1071) );
  inv1f U722 ( .I(n726), .ZN(n1388) );
  inv1f U723 ( .I(n1388), .ZN(n1389) );
  inv1 U725 ( .I(n1388), .ZN(n1390) );
  and2f U731 ( .A1(n1390), .A2(n1071), .Z(n800) );
  and2f U732 ( .A1(n1099), .A2(a), .Z(n719) );
  inv1 U733 ( .I(n1099), .ZN(n726) );
  or2f U734 ( .A1(n1205), .A2(n1362), .Z(n740) );
  inv1f U737 ( .I(i), .ZN(n1362) );
  and2 U738 ( .A1(n), .A2(n728), .Z(n727) );
  inv1 U739 ( .I(a), .ZN(n711) );
  inv1 U741 ( .I(n723), .ZN(n940) );
  and2 U742 ( .A1(n974), .A2(n1391), .Z(n882) );
  and2 U748 ( .A1(n729), .A2(n1261), .Z(n1262) );
  or2 U772 ( .A1(n1169), .A2(n1168), .Z(n1265) );
  or2 U791 ( .A1(n821), .A2(n820), .Z(n825) );
  and2 U806 ( .A1(n1148), .A2(n1122), .Z(n1108) );
  or2 U830 ( .A1(n1216), .A2(n714), .Z(n712) );
  or2 U833 ( .A1(n1217), .A2(n1328), .Z(n714) );
  inv1 U834 ( .I(n1086), .ZN(n1394) );
  or2f U835 ( .A1(n883), .A2(n882), .Z(n721) );
  and2f U837 ( .A1(n1358), .A2(n1252), .Z(n1254) );
  inv1f U852 ( .I(n1358), .ZN(n1370) );
  or2f U856 ( .A1(n983), .A2(n982), .Z(n1358) );
  and2f U859 ( .A1(n780), .A2(n1389), .Z(n781) );
  inv1f U860 ( .I(n1273), .ZN(n1391) );
  inv1f U869 ( .I(n1391), .ZN(n1392) );
  inv1 U880 ( .I(n1391), .ZN(n1393) );
  or2f U881 ( .A1(n1032), .A2(n776), .Z(n779) );
  and2f U882 ( .A1(n1362), .A2(n965), .Z(n968) );
  inv1 U884 ( .I(n1359), .ZN(n1252) );
  or2 U885 ( .A1(n1370), .A2(n1246), .Z(n1245) );
  inv1 U913 ( .I(n850), .ZN(n1063) );
  and2 U918 ( .A1(n1180), .A2(n1249), .Z(n1181) );
  and2 U920 ( .A1(n1317), .A2(n1170), .Z(n1172) );
  or2 U924 ( .A1(n703), .A2(n1196), .Z(n1200) );
  and2 U925 ( .A1(n1082), .A2(n1081), .Z(n1083) );
  inv1 U928 ( .I(n1093), .ZN(n1178) );
  and2 U930 ( .A1(n860), .A2(n859), .Z(n861) );
  and2 U934 ( .A1(n817), .A2(n816), .Z(n818) );
  or2 U935 ( .A1(n1107), .A2(n1106), .Z(n1122) );
  or2 U940 ( .A1(n1105), .A2(n1104), .Z(n1106) );
  or2 U945 ( .A1(n981), .A2(n980), .Z(n982) );
  inv1 U951 ( .I(f), .ZN(n1025) );
  inv1 U961 ( .I(n1122), .ZN(n1149) );
  or2 U962 ( .A1(n823), .A2(m), .Z(n1148) );
  or2 U984 ( .A1(n1282), .A2(n1281), .Z(n1325) );
  or2 U985 ( .A1(n1263), .A2(n1262), .Z(n1282) );
  and2 U986 ( .A1(n1317), .A2(n703), .Z(n1266) );
  and2 U987 ( .A1(n1220), .A2(n1219), .Z(n1221) );
  and2 U993 ( .A1(n1356), .A2(n1355), .Z(n1357) );
  or2f U1002 ( .A1(n1327), .A2(n1326), .Z(n1343) );
  inv1 U1006 ( .I(n1217), .ZN(n1326) );
  or2f U1008 ( .A1(n1249), .A2(n921), .Z(n922) );
  inv1 U1010 ( .I(n912), .ZN(n702) );
  or2f U1011 ( .A1(n1223), .A2(n1222), .Z(n1224) );
  or2f U1013 ( .A1(n1295), .A2(n62), .Z(n1323) );
  and2 U1016 ( .A1(n701), .A2(n1265), .Z(n1171) );
  inv1 U1017 ( .I(n701), .ZN(n1317) );
  and2f U1059 ( .A1(n723), .A2(n1141), .Z(n893) );
  or2f U1063 ( .A1(n1225), .A2(n1224), .Z(q) );
  inv1f U1064 ( .I(n1185), .ZN(n1183) );
  or2f U1067 ( .A1(n1087), .A2(f), .Z(n891) );
  and2f U1075 ( .A1(n1289), .A2(n1288), .Z(n1294) );
  or2f U1076 ( .A1(n993), .A2(n992), .Z(n1284) );
  and2f U1079 ( .A1(n1226), .A2(n1370), .Z(n993) );
  and2f U1081 ( .A1(n711), .A2(e), .Z(n710) );
  or2f U1089 ( .A1(n806), .A2(n805), .Z(n817) );
  inv1 U1090 ( .I(n1071), .ZN(n1078) );
  or2f U1092 ( .A1(n1341), .A2(n1340), .Z(n1354) );
  and2f U1168 ( .A1(n1272), .A2(n1177), .Z(n1193) );
  or2f U1175 ( .A1(n1176), .A2(n1175), .Z(n1177) );
  or2f U1179 ( .A1(n725), .A2(n856), .Z(n860) );
  and2f U1181 ( .A1(n855), .A2(n854), .Z(n856) );
  or2f U1182 ( .A1(n852), .A2(n1064), .Z(n855) );
  inv1f U1191 ( .I(n721), .ZN(n724) );
  or2f U1192 ( .A1(n1260), .A2(n1259), .Z(n1261) );
  or2f U1198 ( .A1(n1179), .A2(n1178), .Z(n1250) );
  or2f U1199 ( .A1(n1251), .A2(n1250), .Z(n1359) );
  or2f U1200 ( .A1(n1221), .A2(n1349), .Z(n1222) );
  and2f U1213 ( .A1(n901), .A2(n900), .Z(n904) );
  and2f U1236 ( .A1(n729), .A2(n1191), .Z(n1192) );
  or2f U1255 ( .A1(n892), .A2(n1063), .Z(n959) );
  or2f U1256 ( .A1(n1213), .A2(n1212), .Z(n1214) );
  and2f U1258 ( .A1(n1226), .A2(n1196), .Z(n987) );
  and2f U1259 ( .A1(n1371), .A2(k), .Z(n723) );
  and2f U1260 ( .A1(n729), .A2(n1098), .Z(n1103) );
  or2f U1264 ( .A1(n1097), .A2(n1096), .Z(n1098) );
  or2f U1265 ( .A1(n1078), .A2(n1390), .Z(n1080) );
  and2f U1267 ( .A1(c), .A2(n1249), .Z(n1251) );
  or2f U1268 ( .A1(n701), .A2(n973), .Z(n915) );
  and2f U1269 ( .A1(n710), .A2(n891), .Z(n892) );
  or2f U1271 ( .A1(l), .A2(n925), .Z(n394) );
  and2f U1279 ( .A1(n1246), .A2(n924), .Z(n925) );
  and2f U1280 ( .A1(n918), .A2(n917), .Z(n920) );
  or2f U1281 ( .A1(n1317), .A2(n974), .Z(n918) );
  or2f U1282 ( .A1(n1326), .A2(n1327), .Z(n1218) );
  or2f U1294 ( .A1(n1193), .A2(n1192), .Z(n1194) );
  and2f U1295 ( .A1(c), .A2(n1196), .Z(n1182) );
  or2f U1296 ( .A1(n893), .A2(n959), .Z(n894) );
  or2f U1297 ( .A1(n1339), .A2(n1338), .Z(n1340) );
  and2f U1298 ( .A1(n1356), .A2(n1343), .Z(n1329) );
  inv1f U1299 ( .I(n1333), .ZN(n1335) );
  or2f U1300 ( .A1(n972), .A2(n971), .Z(n1333) );
  or2f U1301 ( .A1(n970), .A2(n969), .Z(n971) );
  or2f U1322 ( .A1(n819), .A2(n818), .Z(n820) );
  or2f U1327 ( .A1(n1149), .A2(n1148), .Z(n1327) );
  or2f U1328 ( .A1(n822), .A2(n1328), .Z(n823) );
  and2f U1329 ( .A1(n1226), .A2(n1086), .Z(n796) );
  or2f U1330 ( .A1(n760), .A2(n759), .Z(n1099) );
  or2f U1337 ( .A1(n752), .A2(n751), .Z(n760) );
  and2f U1338 ( .A1(n784), .A2(n783), .Z(n1086) );
  and2f U1339 ( .A1(n779), .A2(n778), .Z(n784) );
  and2f U1340 ( .A1(n712), .A2(n713), .Z(n1219) );
  or2f U1355 ( .A1(n1172), .A2(n1171), .Z(n1174) );
  or2f U1360 ( .A1(n1215), .A2(n1214), .Z(n1217) );
  or2f U1364 ( .A1(n1195), .A2(n1194), .Z(n1215) );
  or2f U1384 ( .A1(b), .A2(n1025), .Z(n850) );
  and2f U1385 ( .A1(n1393), .A2(n1197), .Z(n1169) );
  or2f U1386 ( .A1(n873), .A2(n872), .Z(n1273) );
  or2f U1387 ( .A1(n867), .A2(n866), .Z(n873) );
  and2f U1388 ( .A1(n1331), .A2(n1330), .Z(n1339) );
  or2f U1389 ( .A1(n1329), .A2(n1328), .Z(n1330) );
  inv1f U1393 ( .I(n703), .ZN(n709) );
  or2f U1394 ( .A1(n987), .A2(n986), .Z(n703) );
  or2f U1404 ( .A1(n1325), .A2(n1324), .Z(n1356) );
  or2f U1419 ( .A1(n1323), .A2(n1322), .Z(n1324) );
  inv1f U1420 ( .I(n1249), .ZN(n1196) );
  or2f U1421 ( .A1(n920), .A2(n919), .Z(n1249) );
  inv1f U1422 ( .I(b), .ZN(n1087) );
  and2f U1423 ( .A1(n704), .A2(n702), .Z(n701) );
endmodule

