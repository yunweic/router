
module comp ( f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, 
        l, k, j, i, h, g, f, e, d, c, b, a, i0, h0, g0 );
  input f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n, m, l, k,
         j, i, h, g, f, e, d, c, b, a;
  output i0, h0, g0;
  wire   n133, n27, n29, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n119, n120, n121, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151;
  assign i0 = n133;

  and2f U2 ( .A1(n27), .A2(n146), .Z(g0) );
  and2f U7 ( .A1(n35), .A2(n36), .Z(n34) );
  or2f U8 ( .A1(n38), .A2(n37), .Z(n36) );
  and2f U9 ( .A1(n39), .A2(n40), .Z(n38) );
  or2f U11 ( .A1(n42), .A2(n43), .Z(n27) );
  or2f U12 ( .A1(n44), .A2(n45), .Z(n43) );
  or2f U14 ( .A1(n46), .A2(n47), .Z(n40) );
  and2f U15 ( .A1(n48), .A2(n49), .Z(n47) );
  or2f U16 ( .A1(n50), .A2(n51), .Z(n48) );
  and2f U17 ( .A1(n52), .A2(n53), .Z(n51) );
  and2f U19 ( .A1(n55), .A2(n56), .Z(n54) );
  or2f U20 ( .A1(n57), .A2(n58), .Z(n56) );
  or2f U21 ( .A1(n59), .A2(f0), .Z(n57) );
  and2f U30 ( .A1(n69), .A2(n70), .Z(n68) );
  or2f U31 ( .A1(n71), .A2(n72), .Z(n69) );
  or2f U33 ( .A1(n75), .A2(n76), .Z(n73) );
  and2f U35 ( .A1(n78), .A2(n79), .Z(n77) );
  inv1f U49 ( .I(n85), .ZN(n44) );
  and2f U50 ( .A1(n39), .A2(n35), .Z(n85) );
  and2f U51 ( .A1(n86), .A2(n87), .Z(n35) );
  and2f U52 ( .A1(n88), .A2(n89), .Z(n87) );
  inv1f U54 ( .I(n33), .ZN(n88) );
  or2f U55 ( .A1(n91), .A2(n92), .Z(n33) );
  and2f U56 ( .A1(n93), .A2(n94), .Z(n92) );
  or2f U57 ( .A1(n95), .A2(n96), .Z(n93) );
  and2f U58 ( .A1(n97), .A2(n98), .Z(n96) );
  or2f U59 ( .A1(n99), .A2(n100), .Z(n97) );
  and2f U60 ( .A1(n101), .A2(h), .Z(n100) );
  and2f U61 ( .A1(n102), .A2(n90), .Z(n101) );
  or2f U72 ( .A1(g), .A2(n103), .Z(n102) );
  inv1f U73 ( .I(w), .ZN(n103) );
  and2f U74 ( .A1(n107), .A2(n108), .Z(n39) );
  and2f U75 ( .A1(n109), .A2(n110), .Z(n108) );
  inv1f U77 ( .I(n37), .ZN(n109) );
  or2f U78 ( .A1(n113), .A2(n112), .Z(n37) );
  and2f U79 ( .A1(n114), .A2(n115), .Z(n113) );
  and2f U86 ( .A1(k), .A2(n124), .Z(n120) );
  or2f U91 ( .A1(j), .A2(n125), .Z(n119) );
  and2f U101 ( .A1(n60), .A2(e0), .Z(n59) );
  inv1f U109 ( .I(o), .ZN(n60) );
  and2f U110 ( .A1(n77), .A2(d), .Z(n76) );
  or2 U111 ( .A1(n135), .A2(n64), .Z(n45) );
  inv1 U112 ( .I(n150), .ZN(n148) );
  or2 U113 ( .A1(n29), .A2(n136), .Z(n150) );
  and2f U114 ( .A1(n73), .A2(n74), .Z(n72) );
  and2f U115 ( .A1(n83), .A2(n138), .Z(n136) );
  and2f U116 ( .A1(n139), .A2(n140), .Z(n138) );
  inv1 U117 ( .I(b0), .ZN(n111) );
  inv1 U118 ( .I(s), .ZN(n80) );
  inv1 U119 ( .I(x), .ZN(n90) );
  inv1 U120 ( .I(a0), .ZN(n124) );
  inv1 U121 ( .I(n54), .ZN(n52) );
  inv1 U122 ( .I(n137), .ZN(n139) );
  inv1 U123 ( .I(n68), .ZN(n140) );
  or2 U124 ( .A1(n67), .A2(n68), .Z(n29) );
  inv1 U125 ( .I(z), .ZN(n134) );
  inv1 U126 ( .I(z), .ZN(n125) );
  or2 U127 ( .A1(n63), .A2(n40), .Z(n135) );
  or2 U128 ( .A1(n67), .A2(n65), .Z(n137) );
  inv1 U129 ( .I(n138), .ZN(n64) );
  and2f U130 ( .A1(j), .A2(n134), .Z(n116) );
  or2f U131 ( .A1(n124), .A2(k), .Z(n141) );
  and2f U132 ( .A1(n141), .A2(n142), .Z(n121) );
  and2f U133 ( .A1(l), .A2(n111), .Z(n142) );
  or2f U134 ( .A1(n121), .A2(n145), .Z(n143) );
  and2f U135 ( .A1(n143), .A2(n144), .Z(n114) );
  or2 U136 ( .A1(n116), .A2(n119), .Z(n144) );
  or2f U137 ( .A1(n120), .A2(n116), .Z(n145) );
  or2 U138 ( .A1(k), .A2(n124), .Z(n123) );
  or2f U139 ( .A1(n147), .A2(n148), .Z(n146) );
  inv1 U140 ( .I(n146), .ZN(n133) );
  inv1f U141 ( .I(n149), .ZN(n147) );
  or2f U142 ( .A1(n34), .A2(n151), .Z(n149) );
  or2 U143 ( .A1(n33), .A2(n29), .Z(n151) );
  or2 U144 ( .A1(f), .A2(n104), .Z(n98) );
  inv1 U145 ( .I(v), .ZN(n104) );
  or2 U146 ( .A1(b), .A2(n81), .Z(n74) );
  inv1 U147 ( .I(d0), .ZN(n61) );
  inv1 U148 ( .I(y), .ZN(n126) );
  or2 U149 ( .A1(i), .A2(n126), .Z(n115) );
  and2 U150 ( .A1(n102), .A2(n106), .Z(n86) );
  and2 U151 ( .A1(n94), .A2(n98), .Z(n106) );
  and2 U152 ( .A1(a), .A2(n82), .Z(n67) );
  inv1 U153 ( .I(t), .ZN(n79) );
  inv1 U154 ( .I(r), .ZN(n81) );
  or2 U155 ( .A1(n111), .A2(l), .Z(n110) );
  inv1 U156 ( .I(p), .ZN(n58) );
  and2 U157 ( .A1(i), .A2(n126), .Z(n112) );
  and2 U158 ( .A1(m), .A2(n62), .Z(n46) );
  and2 U159 ( .A1(f0), .A2(n58), .Z(n130) );
  inv1 U160 ( .I(n131), .ZN(n128) );
  and2 U161 ( .A1(n49), .A2(n53), .Z(n131) );
  and2 U162 ( .A1(e), .A2(n105), .Z(n91) );
  inv1 U163 ( .I(n83), .ZN(n63) );
  and2 U164 ( .A1(n78), .A2(n84), .Z(n83) );
  or2 U165 ( .A1(n60), .A2(e0), .Z(n55) );
  and2 U166 ( .A1(n), .A2(n61), .Z(n50) );
  inv1 U167 ( .I(c0), .ZN(n62) );
  or2 U168 ( .A1(n90), .A2(h), .Z(n89) );
  or2 U169 ( .A1(n), .A2(n61), .Z(n53) );
  or2 U170 ( .A1(m), .A2(n62), .Z(n49) );
  and2 U171 ( .A1(c), .A2(n80), .Z(n75) );
  and2 U172 ( .A1(b), .A2(n81), .Z(n71) );
  inv1 U173 ( .I(q), .ZN(n82) );
  or2 U174 ( .A1(a), .A2(n82), .Z(n70) );
  and2 U175 ( .A1(n123), .A2(n127), .Z(n107) );
  and2 U176 ( .A1(n115), .A2(n119), .Z(n127) );
  inv1 U177 ( .I(u), .ZN(n105) );
  or2 U178 ( .A1(e), .A2(n105), .Z(n94) );
  and2 U179 ( .A1(g), .A2(n103), .Z(n99) );
  and2 U180 ( .A1(f), .A2(n104), .Z(n95) );
  or2 U181 ( .A1(c), .A2(n80), .Z(n78) );
  and2 U182 ( .A1(n70), .A2(n74), .Z(n84) );
  and2 U183 ( .A1(t), .A2(n66), .Z(n65) );
  inv1 U184 ( .I(d), .ZN(n66) );
  or2 U185 ( .A1(n128), .A2(n129), .Z(n42) );
  or2 U186 ( .A1(n59), .A2(n130), .Z(n129) );
  inv1 U187 ( .I(n27), .ZN(h0) );
endmodule

