
module x1 ( z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, 
        i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, w, v, u, t, s, r, q, p, o, n, 
        m, l, k, j, i, h, g, f, e, d, c, b, a, i2, h2, g2, f2, e2, d2, c2, b2, 
        a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, 
        i1, h1, g1, f1, e1, d1, c1, b1, a1 );
  input z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0,
         h0, g0, f0, e0, d0, c0, b0, a0, z, y, w, v, u, t, s, r, q, p, o, n, m,
         l, k, j, i, h, g, f, e, d, c, b, a;
  output i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1,
         r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1,
         a1;
  wire   n341, n342, n343, n344, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n345, n346, n347, n348, n349;

  and2f U51 ( .A1(n106), .A2(n107), .Z(n96) );
  and2f U52 ( .A1(n108), .A2(n109), .Z(n106) );
  or2f U53 ( .A1(n110), .A2(n111), .Z(n108) );
  or2f U59 ( .A1(n116), .A2(n117), .Z(n110) );
  or2f U74 ( .A1(n138), .A2(n139), .Z(l1) );
  or2f U75 ( .A1(n140), .A2(n141), .Z(n139) );
  and2f U77 ( .A1(n142), .A2(n143), .Z(n140) );
  or2f U78 ( .A1(n144), .A2(n145), .Z(n142) );
  and2f U83 ( .A1(o), .A2(n151), .Z(n148) );
  or2f U84 ( .A1(n152), .A2(n153), .Z(n151) );
  or2f U86 ( .A1(n137), .A2(e0), .Z(n150) );
  and2f U88 ( .A1(p), .A2(n126), .Z(n154) );
  or2f U102 ( .A1(n45), .A2(n168), .Z(n167) );
  or2f U138 ( .A1(n205), .A2(n206), .Z(n200) );
  or2f U156 ( .A1(n221), .A2(n222), .Z(g2) );
  or2f U157 ( .A1(n223), .A2(n224), .Z(n222) );
  or2f U165 ( .A1(n232), .A2(v), .Z(n231) );
  and2f U166 ( .A1(o), .A2(n233), .Z(n232) );
  or2f U167 ( .A1(n234), .A2(n235), .Z(n233) );
  and2f U171 ( .A1(n238), .A2(n239), .Z(n229) );
  and2f U177 ( .A1(n241), .A2(p0), .Z(n238) );
  and2f U182 ( .A1(n123), .A2(n247), .Z(n246) );
  or2f U183 ( .A1(n103), .A2(n248), .Z(n123) );
  and2f U191 ( .A1(n253), .A2(a0), .Z(n225) );
  and2f U193 ( .A1(n255), .A2(l), .Z(n254) );
  and2f U194 ( .A1(b), .A2(n256), .Z(n255) );
  and2f U227 ( .A1(d), .A2(d0), .Z(n137) );
  and2f U239 ( .A1(n291), .A2(i), .Z(n290) );
  and2f U240 ( .A1(n292), .A2(n349), .Z(n291) );
  and2f U244 ( .A1(n278), .A2(n92), .Z(n294) );
  or2f U245 ( .A1(n265), .A2(n130), .Z(n92) );
  or2f U246 ( .A1(n285), .A2(n127), .Z(n265) );
  and2f U249 ( .A1(q0), .A2(n81), .Z(n295) );
  or2f U256 ( .A1(n285), .A2(n130), .Z(n268) );
  and2f U258 ( .A1(n81), .A2(n349), .Z(n53) );
  inv1f U274 ( .I(p), .ZN(n130) );
  or2f U279 ( .A1(e), .A2(u), .Z(n143) );
  and2f U290 ( .A1(n82), .A2(n314), .Z(n203) );
  and2f U292 ( .A1(l), .A2(n316), .Z(n82) );
  and2f U293 ( .A1(n349), .A2(b), .Z(n316) );
  buf0 U319 ( .I(m0), .Z(i1) );
  buf0 U320 ( .I(n0), .Z(j1) );
  buf0 U321 ( .I(y), .Z(p1) );
  buf0 U322 ( .I(z), .Z(q1) );
  buf0 U323 ( .I(n344), .Z(s1) );
  buf0 U324 ( .I(x0), .Z(t1) );
  buf0 U325 ( .I(y0), .Z(u1) );
  buf0 U326 ( .I(n343), .Z(x1) );
  buf0 U327 ( .I(n342), .Z(z1) );
  buf0 U328 ( .I(n341), .Z(a2) );
  buf0 U329 ( .I(h0), .Z(c2) );
  or2 U330 ( .A1(n196), .A2(n194), .Z(n205) );
  and2f U331 ( .A1(n203), .A2(n207), .Z(n194) );
  and2f U332 ( .A1(a0), .A2(n203), .Z(n196) );
  and2 U333 ( .A1(n107), .A2(p), .Z(n235) );
  and2f U334 ( .A1(n247), .A2(n305), .Z(n107) );
  and2 U335 ( .A1(n154), .A2(d0), .Z(n152) );
  or2 U336 ( .A1(v), .A2(g), .Z(n245) );
  inv1 U337 ( .I(n254), .ZN(n253) );
  and2 U338 ( .A1(n246), .A2(n121), .Z(n243) );
  and2 U339 ( .A1(n150), .A2(n126), .Z(n149) );
  inv1 U340 ( .I(g), .ZN(n126) );
  and2 U341 ( .A1(n284), .A2(n285), .Z(n283) );
  or2 U342 ( .A1(n286), .A2(n287), .Z(n284) );
  and2 U343 ( .A1(a), .A2(n165), .Z(n163) );
  or2 U344 ( .A1(n166), .A2(n167), .Z(n165) );
  or2 U345 ( .A1(n183), .A2(n184), .Z(n182) );
  or2 U346 ( .A1(n185), .A2(n169), .Z(n184) );
  or2 U347 ( .A1(n112), .A2(n113), .Z(n111) );
  inv1 U348 ( .I(n345), .ZN(n46) );
  or2 U349 ( .A1(n293), .A2(n88), .Z(n292) );
  and2 U350 ( .A1(n294), .A2(g), .Z(n293) );
  or2 U351 ( .A1(n229), .A2(n230), .Z(n228) );
  and2 U352 ( .A1(d0), .A2(n231), .Z(n230) );
  or2 U353 ( .A1(n252), .A2(n225), .Z(n250) );
  or2 U354 ( .A1(n344), .A2(n226), .Z(n221) );
  or2 U355 ( .A1(n193), .A2(n199), .Z(n198) );
  and2 U356 ( .A1(n200), .A2(n201), .Z(n199) );
  and2f U357 ( .A1(n73), .A2(n74), .Z(n72) );
  and2 U358 ( .A1(h), .A2(n220), .Z(n223) );
  or2 U359 ( .A1(m), .A2(j), .Z(n345) );
  inv1 U360 ( .I(m), .ZN(n247) );
  inv1 U361 ( .I(j), .ZN(n42) );
  inv1f U362 ( .I(n123), .ZN(n122) );
  inv1 U363 ( .I(v), .ZN(n81) );
  or2f U364 ( .A1(n295), .A2(p0), .Z(n278) );
  and2f U365 ( .A1(q0), .A2(n128), .Z(n124) );
  inv1 U366 ( .I(n268), .ZN(n128) );
  inv1 U367 ( .I(n143), .ZN(n305) );
  or2 U368 ( .A1(n71), .A2(z0), .Z(n256) );
  and2f U369 ( .A1(n46), .A2(r), .Z(n71) );
  or2f U370 ( .A1(n148), .A2(n348), .Z(n346) );
  and2 U371 ( .A1(n346), .A2(n347), .Z(n145) );
  or2 U372 ( .A1(h0), .A2(n53), .Z(n347) );
  or2 U373 ( .A1(n149), .A2(h0), .Z(n348) );
  and2f U374 ( .A1(n120), .A2(n121), .Z(n119) );
  or2f U375 ( .A1(n63), .A2(n64), .Z(n62) );
  and2f U376 ( .A1(n71), .A2(n72), .Z(n63) );
  and2f U377 ( .A1(n150), .A2(n130), .Z(n153) );
  or2f U378 ( .A1(n118), .A2(n119), .Z(n117) );
  and2f U379 ( .A1(n124), .A2(n125), .Z(n118) );
  or2f U380 ( .A1(n75), .A2(n76), .Z(n73) );
  and2f U381 ( .A1(n78), .A2(n79), .Z(n75) );
  inv1f U382 ( .I(a), .ZN(n349) );
  inv1 U383 ( .I(w), .ZN(n109) );
  and2 U384 ( .A1(n315), .A2(n247), .Z(n314) );
  inv1 U385 ( .I(n92), .ZN(n158) );
  and2 U386 ( .A1(n247), .A2(n67), .Z(n101) );
  or2 U387 ( .A1(n126), .A2(n68), .Z(n94) );
  or2 U388 ( .A1(p0), .A2(q0), .Z(n91) );
  and2 U389 ( .A1(n248), .A2(d0), .Z(n260) );
  and2 U390 ( .A1(n285), .A2(e0), .Z(n261) );
  or2 U391 ( .A1(j), .A2(v), .Z(n197) );
  and2 U392 ( .A1(g0), .A2(j), .Z(n102) );
  or2 U393 ( .A1(n324), .A2(n325), .Z(n323) );
  or2 U394 ( .A1(n322), .A2(n326), .Z(n325) );
  or2 U395 ( .A1(n327), .A2(n328), .Z(n324) );
  inv1 U396 ( .I(l), .ZN(n326) );
  inv1 U397 ( .I(b), .ZN(n322) );
  and2 U398 ( .A1(n313), .A2(n196), .Z(n312) );
  and2 U399 ( .A1(n197), .A2(n80), .Z(n313) );
  and2 U400 ( .A1(n317), .A2(n318), .Z(n311) );
  and2 U401 ( .A1(b), .A2(n46), .Z(n317) );
  and2 U402 ( .A1(n319), .A2(n56), .Z(n318) );
  and2 U403 ( .A1(n349), .A2(n315), .Z(n319) );
  and2 U404 ( .A1(n310), .A2(c), .Z(n308) );
  and2 U405 ( .A1(n102), .A2(n109), .Z(n310) );
  and2 U406 ( .A1(t0), .A2(o0), .Z(n309) );
  and2 U407 ( .A1(n53), .A2(n268), .Z(n301) );
  and2 U408 ( .A1(n260), .A2(n101), .Z(n300) );
  or2 U409 ( .A1(v), .A2(n247), .Z(n299) );
  and2 U410 ( .A1(n283), .A2(n137), .Z(n282) );
  and2 U411 ( .A1(n288), .A2(g), .Z(n286) );
  and2 U412 ( .A1(n267), .A2(n261), .Z(n281) );
  and2 U413 ( .A1(n101), .A2(n349), .Z(n267) );
  and2 U414 ( .A1(e0), .A2(n128), .Z(n266) );
  and2 U415 ( .A1(n94), .A2(n265), .Z(n264) );
  and2 U416 ( .A1(n240), .A2(n180), .Z(n239) );
  and2 U417 ( .A1(n349), .A2(n67), .Z(n240) );
  and2 U418 ( .A1(n220), .A2(n349), .Z(n219) );
  or2 U419 ( .A1(n218), .A2(e), .Z(n217) );
  or2 U420 ( .A1(u), .A2(w), .Z(n218) );
  or2 U421 ( .A1(n171), .A2(n172), .Z(n166) );
  and2 U422 ( .A1(r0), .A2(b), .Z(n164) );
  and2 U423 ( .A1(m), .A2(n182), .Z(n175) );
  or2 U424 ( .A1(e0), .A2(n189), .Z(n183) );
  or2 U425 ( .A1(n177), .A2(n178), .Z(n176) );
  and2 U426 ( .A1(n44), .A2(n179), .Z(n178) );
  and2 U427 ( .A1(n181), .A2(w), .Z(n177) );
  or2 U428 ( .A1(l0), .A2(p0), .Z(n179) );
  or2 U429 ( .A1(n160), .A2(f0), .Z(n159) );
  and2 U430 ( .A1(k), .A2(a0), .Z(n160) );
  and2 U431 ( .A1(h), .A2(n155), .Z(n144) );
  and2 U432 ( .A1(w), .A2(h0), .Z(n141) );
  and2 U433 ( .A1(n158), .A2(n91), .Z(n157) );
  and2 U434 ( .A1(n136), .A2(n137), .Z(n133) );
  and2 U435 ( .A1(n135), .A2(n130), .Z(n134) );
  and2 U436 ( .A1(n100), .A2(n101), .Z(n99) );
  and2 U437 ( .A1(n102), .A2(n103), .Z(n100) );
  and2 U438 ( .A1(n104), .A2(n105), .Z(n98) );
  and2 U439 ( .A1(f), .A2(g0), .Z(n104) );
  and2 U440 ( .A1(v), .A2(n42), .Z(n105) );
  and2 U441 ( .A1(n93), .A2(n53), .Z(n89) );
  inv1 U442 ( .I(n94), .ZN(n93) );
  and2 U443 ( .A1(n91), .A2(n92), .Z(n90) );
  and2 U444 ( .A1(n86), .A2(n349), .Z(n85) );
  or2 U445 ( .A1(n87), .A2(n88), .Z(n86) );
  and2 U446 ( .A1(i0), .A2(n67), .Z(n87) );
  or2 U447 ( .A1(n59), .A2(n53), .Z(n58) );
  and2 U448 ( .A1(n349), .A2(n60), .Z(n59) );
  inv1 U449 ( .I(f), .ZN(n60) );
  or2 U450 ( .A1(n50), .A2(n51), .Z(n49) );
  and2 U451 ( .A1(n55), .A2(n), .Z(n50) );
  and2 U452 ( .A1(n52), .A2(n53), .Z(n51) );
  and2 U453 ( .A1(n56), .A2(n349), .Z(n55) );
  or2 U454 ( .A1(n130), .A2(n126), .Z(n237) );
  and2 U455 ( .A1(n107), .A2(n304), .Z(n136) );
  and2 U456 ( .A1(n349), .A2(o), .Z(n304) );
  or2 U457 ( .A1(e0), .A2(p0), .Z(n170) );
  and2 U458 ( .A1(n81), .A2(n109), .Z(n135) );
  or2 U459 ( .A1(n273), .A2(n274), .Z(n271) );
  or2 U460 ( .A1(n276), .A2(n277), .Z(n273) );
  or2 U461 ( .A1(n275), .A2(n68), .Z(n274) );
  or2 U462 ( .A1(a), .A2(n121), .Z(n277) );
  inv1 U463 ( .I(i0), .ZN(n272) );
  or2 U464 ( .A1(h0), .A2(n296), .Z(n210) );
  or2 U465 ( .A1(z), .A2(y), .Z(n296) );
  and2 U466 ( .A1(n257), .A2(h), .Z(n252) );
  or2 U467 ( .A1(n220), .A2(n173), .Z(n257) );
  or2 U468 ( .A1(f0), .A2(r0), .Z(n341) );
  or2 U469 ( .A1(m0), .A2(x0), .Z(n226) );
  or2 U470 ( .A1(n258), .A2(n259), .Z(n220) );
  or2 U471 ( .A1(s0), .A2(p0), .Z(n258) );
  or2 U472 ( .A1(n260), .A2(n261), .Z(n259) );
  and2 U473 ( .A1(n42), .A2(n56), .Z(n207) );
  and2 U474 ( .A1(n196), .A2(n197), .Z(n195) );
  or2 U475 ( .A1(n208), .A2(n209), .Z(n193) );
  or2 U476 ( .A1(n137), .A2(n214), .Z(n208) );
  or2 U477 ( .A1(n210), .A2(n211), .Z(n209) );
  or2 U478 ( .A1(c0), .A2(b0), .Z(n214) );
  and2 U479 ( .A1(c), .A2(n102), .Z(n192) );
  inv1 U480 ( .I(q), .ZN(n127) );
  and2 U481 ( .A1(n126), .A2(n127), .Z(n125) );
  inv1 U482 ( .I(r), .ZN(n54) );
  inv1 U483 ( .I(d), .ZN(n248) );
  inv1 U484 ( .I(n329), .ZN(n327) );
  or2 U485 ( .A1(n197), .A2(r), .Z(n329) );
  or2 U486 ( .A1(n), .A2(m), .Z(n328) );
  inv1 U487 ( .I(k), .ZN(n80) );
  inv1 U488 ( .I(n), .ZN(n315) );
  inv1 U489 ( .I(o), .ZN(n285) );
  and2 U490 ( .A1(n143), .A2(n247), .Z(n288) );
  and2 U491 ( .A1(n107), .A2(n109), .Z(n287) );
  inv1 U492 ( .I(n236), .ZN(n234) );
  or2 U493 ( .A1(n237), .A2(m), .Z(n236) );
  and2 U494 ( .A1(n242), .A2(n92), .Z(n241) );
  or2 U495 ( .A1(n243), .A2(n244), .Z(n242) );
  and2 U496 ( .A1(n245), .A2(n68), .Z(n244) );
  or2 U497 ( .A1(n169), .A2(n170), .Z(n168) );
  or2 U498 ( .A1(n173), .A2(n174), .Z(n172) );
  and2 U499 ( .A1(g0), .A2(n42), .Z(n174) );
  or2 U500 ( .A1(j0), .A2(d0), .Z(n171) );
  or2 U501 ( .A1(h0), .A2(n186), .Z(n169) );
  or2 U502 ( .A1(s0), .A2(q0), .Z(n186) );
  and2 U503 ( .A1(n187), .A2(n81), .Z(n185) );
  or2 U504 ( .A1(n342), .A2(n188), .Z(n187) );
  or2 U505 ( .A1(p0), .A2(b0), .Z(n188) );
  or2 U506 ( .A1(k0), .A2(g0), .Z(n189) );
  and2 U507 ( .A1(n137), .A2(n81), .Z(n181) );
  or2 U508 ( .A1(d0), .A2(e0), .Z(n155) );
  and2 U509 ( .A1(n122), .A2(p0), .Z(n120) );
  and2 U510 ( .A1(n129), .A2(e0), .Z(n116) );
  and2 U511 ( .A1(o), .A2(n130), .Z(n129) );
  or2 U512 ( .A1(n114), .A2(n115), .Z(n113) );
  and2 U513 ( .A1(s0), .A2(n67), .Z(n114) );
  and2 U514 ( .A1(h0), .A2(n42), .Z(n115) );
  and2 U515 ( .A1(w0), .A2(o0), .Z(n112) );
  inv1 U516 ( .I(c), .ZN(n103) );
  inv1 U517 ( .I(h), .ZN(n67) );
  inv1 U518 ( .I(s), .ZN(n74) );
  and2 U519 ( .A1(n53), .A2(k0), .Z(n77) );
  and2 U520 ( .A1(n80), .A2(n81), .Z(n79) );
  and2 U521 ( .A1(a0), .A2(n82), .Z(n78) );
  and2 U522 ( .A1(k0), .A2(n54), .Z(n52) );
  or2 U523 ( .A1(n54), .A2(n74), .Z(n180) );
  and2 U524 ( .A1(p0), .A2(v), .Z(n88) );
  inv1 U525 ( .I(n245), .ZN(n121) );
  and2 U526 ( .A1(n158), .A2(n81), .Z(n275) );
  inv1 U527 ( .I(n278), .ZN(n276) );
  inv1 U528 ( .I(i), .ZN(n68) );
  and2 U529 ( .A1(i0), .A2(t), .Z(n173) );
  and2 U530 ( .A1(k0), .A2(v), .Z(n56) );
  or2 U531 ( .A1(n212), .A2(n213), .Z(n211) );
  and2 U532 ( .A1(i), .A2(i0), .Z(n213) );
  and2 U533 ( .A1(d0), .A2(n67), .Z(n212) );
  and2 U534 ( .A1(i0), .A2(n69), .Z(n65) );
  inv1 U535 ( .I(n70), .ZN(n69) );
  and2 U536 ( .A1(t), .A2(a), .Z(n70) );
  and2 U537 ( .A1(n67), .A2(n68), .Z(n66) );
  and2 U538 ( .A1(n77), .A2(b), .Z(n76) );
  or2 U539 ( .A1(a0), .A2(k0), .Z(n45) );
  inv1 U540 ( .I(n180), .ZN(n44) );
  or2 U541 ( .A1(n40), .A2(n41), .Z(n343) );
  or2 U542 ( .A1(z), .A2(h0), .Z(n41) );
  and2 U543 ( .A1(n42), .A2(n43), .Z(n40) );
  or2 U544 ( .A1(g0), .A2(n341), .Z(n43) );
  or2 U545 ( .A1(c0), .A2(d0), .Z(n342) );
  or2 U546 ( .A1(n341), .A2(n225), .Z(n224) );
  and2 U547 ( .A1(n173), .A2(h), .Z(n344) );
  and2 U548 ( .A1(g0), .A2(c), .Z(n206) );
  or2 U549 ( .A1(j), .A2(n202), .Z(n201) );
  and2 U550 ( .A1(n203), .A2(n204), .Z(n202) );
  and2 U551 ( .A1(n45), .A2(v), .Z(n204) );
  and2 U552 ( .A1(n341), .A2(n322), .Z(n321) );
  and2 U553 ( .A1(a0), .A2(n323), .Z(n320) );
  or2 U554 ( .A1(n308), .A2(n309), .Z(n307) );
  or2 U555 ( .A1(n311), .A2(n312), .Z(n306) );
  and2 U556 ( .A1(c0), .A2(n299), .Z(n298) );
  and2 U557 ( .A1(n300), .A2(n301), .Z(n297) );
  and2 U558 ( .A1(u0), .A2(o0), .Z(n279) );
  or2 U559 ( .A1(n281), .A2(n282), .Z(n280) );
  and2 U560 ( .A1(n264), .A2(q0), .Z(n263) );
  and2 U561 ( .A1(n266), .A2(n267), .Z(n262) );
  and2 U562 ( .A1(v0), .A2(o0), .Z(n227) );
  inv1 U563 ( .I(n217), .ZN(n216) );
  and2 U564 ( .A1(n219), .A2(h), .Z(n215) );
  or2 U565 ( .A1(n175), .A2(n176), .Z(n161) );
  or2 U566 ( .A1(n163), .A2(n164), .Z(n162) );
  or2 U567 ( .A1(n156), .A2(n157), .Z(n138) );
  and2 U568 ( .A1(b), .A2(n159), .Z(n156) );
  and2 U569 ( .A1(h0), .A2(j), .Z(n132) );
  and2 U570 ( .A1(n133), .A2(n134), .Z(n131) );
  and2 U571 ( .A1(n95), .A2(n349), .Z(n1) );
  or2 U572 ( .A1(n96), .A2(n97), .Z(n95) );
  or2 U573 ( .A1(n98), .A2(n99), .Z(n97) );
  and2 U574 ( .A1(n85), .A2(i), .Z(n84) );
  and2 U575 ( .A1(n89), .A2(n90), .Z(n83) );
  or2 U576 ( .A1(n61), .A2(n62), .Z(r1) );
  and2 U577 ( .A1(j0), .A2(n349), .Z(n61) );
  and2 U578 ( .A1(n65), .A2(n66), .Z(n64) );
  or2 U579 ( .A1(n48), .A2(n49), .Z(n47) );
  and2 U580 ( .A1(g0), .A2(n58), .Z(n48) );
  and2 U581 ( .A1(n135), .A2(n170), .Z(n303) );
  and2 U582 ( .A1(n136), .A2(n237), .Z(n302) );
  or2 U583 ( .A1(i0), .A2(n290), .Z(n289) );
  inv1 U584 ( .I(n210), .ZN(n270) );
  and2 U585 ( .A1(n271), .A2(n272), .Z(n269) );
  or2 U586 ( .A1(n250), .A2(n251), .Z(n249) );
  or2 U587 ( .A1(n226), .A2(n341), .Z(n251) );
  or2 U588 ( .A1(n192), .A2(n193), .Z(n191) );
  or2 U589 ( .A1(n194), .A2(n195), .Z(n190) );
  or2 U590 ( .A1(n320), .A2(n321), .Z(a1) );
  or2 U591 ( .A1(n306), .A2(n307), .Z(b1) );
  and2 U592 ( .A1(b0), .A2(n299), .Z(c1) );
  or2 U593 ( .A1(n297), .A2(n298), .Z(d1) );
  or2 U594 ( .A1(n279), .A2(n280), .Z(e1) );
  or2 U595 ( .A1(n262), .A2(n263), .Z(f1) );
  or2 U596 ( .A1(n227), .A2(n228), .Z(g1) );
  and2 U597 ( .A1(n215), .A2(n216), .Z(h1) );
  or2 U598 ( .A1(n161), .A2(n162), .Z(k1) );
  or2 U599 ( .A1(n131), .A2(n132), .Z(m1) );
  or2 U600 ( .A1(n83), .A2(n84), .Z(o1) );
  and2 U601 ( .A1(n46), .A2(n47), .Z(v1) );
  and2 U602 ( .A1(n44), .A2(n45), .Z(w1) );
  inv1 U603 ( .I(n343), .ZN(y1) );
  and2 U604 ( .A1(n302), .A2(n303), .Z(b2) );
  or2 U605 ( .A1(n210), .A2(n289), .Z(d2) );
  and2 U606 ( .A1(n269), .A2(n270), .Z(e2) );
  inv1 U607 ( .I(n249), .ZN(f2) );
  inv1 U608 ( .I(n198), .ZN(h2) );
  or2 U609 ( .A1(n190), .A2(n191), .Z(i2) );
endmodule

