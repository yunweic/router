
module C432_iscas ( j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, 
        t, s, r, q, p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a, q0, p0, o0, 
        n0, m0, l0, k0 );
  input j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q,
         p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output q0, p0, o0, n0, m0, l0, k0;
  wire   n431, n207, n208, n210, n211, n212, n213, n214, n216, n217, n218,
         n219, n220, n222, n224, n225, n226, n227, n228, n229, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428;

  or2 U215 ( .A1(n287), .A2(n288), .Z(n208) );
  or2 U217 ( .A1(n208), .A2(n212), .Z(n210) );
  or2 U219 ( .A1(n356), .A2(h), .Z(n211) );
  or2 U220 ( .A1(n299), .A2(n356), .Z(n212) );
  or2 U221 ( .A1(w), .A2(n324), .Z(n213) );
  inv1 U222 ( .I(n222), .ZN(n214) );
  or2 U224 ( .A1(n217), .A2(n218), .Z(n216) );
  inv1 U225 ( .I(n359), .ZN(n217) );
  inv1 U226 ( .I(n358), .ZN(n218) );
  or2 U228 ( .A1(o), .A2(n303), .Z(n220) );
  inv1 U231 ( .I(n378), .ZN(l0) );
  and2 U232 ( .A1(n400), .A2(n225), .Z(n224) );
  inv1 U233 ( .I(n403), .ZN(n225) );
  inv1 U235 ( .I(n340), .ZN(n227) );
  and2 U236 ( .A1(n222), .A2(d), .Z(n228) );
  and2 U237 ( .A1(m0), .A2(e), .Z(n229) );
  or2 U240 ( .A1(n311), .A2(n232), .Z(n350) );
  or2 U241 ( .A1(n310), .A2(c), .Z(n232) );
  or2 U243 ( .A1(n316), .A2(a0), .Z(n233) );
  or2 U244 ( .A1(n302), .A2(n234), .Z(n341) );
  or2 U245 ( .A1(n301), .A2(s), .Z(n234) );
  or2 U246 ( .A1(n323), .A2(n235), .Z(n339) );
  or2 U247 ( .A1(n322), .A2(i0), .Z(n235) );
  and2 U248 ( .A1(n238), .A2(n237), .Z(n236) );
  inv1 U249 ( .I(n348), .ZN(n237) );
  inv1 U251 ( .I(n347), .ZN(n239) );
  or2 U254 ( .A1(n236), .A2(n243), .Z(n242) );
  inv1 U255 ( .I(n349), .ZN(n243) );
  or2 U256 ( .A1(n334), .A2(n244), .Z(n338) );
  or2 U257 ( .A1(n401), .A2(i), .Z(n244) );
  or2 U259 ( .A1(n368), .A2(m), .Z(n245) );
  and2 U260 ( .A1(n380), .A2(n381), .Z(n246) );
  or2 U262 ( .A1(n394), .A2(c0), .Z(n247) );
  inv1 U264 ( .I(n248), .ZN(n250) );
  and2 U265 ( .A1(n275), .A2(h), .Z(n249) );
  inv1 U267 ( .I(n385), .ZN(n252) );
  or2 U268 ( .A1(n351), .A2(n253), .Z(n352) );
  or2 U269 ( .A1(n406), .A2(e), .Z(n253) );
  or2 U271 ( .A1(g), .A2(n333), .Z(n255) );
  or2 U275 ( .A1(n363), .A2(u), .Z(n258) );
  inv1 U276 ( .I(d), .ZN(n259) );
  inv1 U278 ( .I(n260), .ZN(n416) );
  inv1 U279 ( .I(n365), .ZN(n261) );
  inv1 U281 ( .I(n388), .ZN(n263) );
  and2 U284 ( .A1(n367), .A2(n277), .Z(n266) );
  or2 U288 ( .A1(n250), .A2(n268), .Z(n270) );
  or2 U293 ( .A1(n208), .A2(n299), .Z(n275) );
  inv1 U295 ( .I(n266), .ZN(n425) );
  inv1 U296 ( .I(n370), .ZN(n277) );
  inv1 U297 ( .I(l), .ZN(n278) );
  and2 U298 ( .A1(n), .A2(n278), .Z(n281) );
  inv1 U299 ( .I(p), .ZN(n279) );
  and2 U300 ( .A1(r), .A2(n279), .Z(n280) );
  or2 U301 ( .A1(n281), .A2(n280), .Z(n288) );
  and2 U302 ( .A1(f), .A2(n259), .Z(n284) );
  inv1 U303 ( .I(a), .ZN(n282) );
  and2 U304 ( .A1(n282), .A2(b), .Z(n283) );
  inv1 U306 ( .I(h), .ZN(n306) );
  and2 U307 ( .A1(j), .A2(n306), .Z(n285) );
  inv1 U310 ( .I(t), .ZN(n289) );
  and2 U311 ( .A1(v), .A2(n289), .Z(n292) );
  inv1 U312 ( .I(x), .ZN(n290) );
  and2 U313 ( .A1(z), .A2(n290), .Z(n291) );
  inv1 U315 ( .I(b0), .ZN(n293) );
  and2 U316 ( .A1(d0), .A2(n293), .Z(n296) );
  inv1 U317 ( .I(f0), .ZN(n294) );
  and2 U318 ( .A1(h0), .A2(n294), .Z(n295) );
  and2 U321 ( .A1(p), .A2(k0), .Z(n302) );
  inv1 U322 ( .I(r), .ZN(n301) );
  or2 U323 ( .A1(n302), .A2(n301), .Z(n363) );
  inv1 U324 ( .I(n341), .ZN(n305) );
  and2 U325 ( .A1(l), .A2(k0), .Z(n304) );
  inv1 U326 ( .I(n), .ZN(n303) );
  or2 U327 ( .A1(n304), .A2(n303), .Z(n372) );
  inv1 U330 ( .I(j), .ZN(n356) );
  inv1 U332 ( .I(n355), .ZN(n309) );
  inv1 U333 ( .I(f), .ZN(n333) );
  or2 U334 ( .A1(n228), .A2(n255), .Z(n332) );
  inv1 U335 ( .I(n332), .ZN(n308) );
  or2 U336 ( .A1(n308), .A2(n309), .Z(n313) );
  and2 U337 ( .A1(a), .A2(k0), .Z(n311) );
  inv1 U338 ( .I(b), .ZN(n310) );
  or2 U339 ( .A1(n311), .A2(n310), .Z(n406) );
  inv1 U340 ( .I(n350), .ZN(n312) );
  and2 U343 ( .A1(x), .A2(k0), .Z(n317) );
  inv1 U344 ( .I(z), .ZN(n316) );
  or2 U345 ( .A1(n317), .A2(n316), .Z(n394) );
  inv1 U346 ( .I(n335), .ZN(n321) );
  inv1 U348 ( .I(d0), .ZN(n318) );
  or2 U350 ( .A1(n390), .A2(e0), .Z(n344) );
  inv1 U351 ( .I(n344), .ZN(n320) );
  or2 U352 ( .A1(n321), .A2(n320), .Z(n329) );
  inv1 U354 ( .I(h0), .ZN(n322) );
  or2 U355 ( .A1(n323), .A2(n322), .Z(n376) );
  inv1 U356 ( .I(n339), .ZN(n327) );
  and2 U357 ( .A1(k0), .A2(t), .Z(n325) );
  inv1 U358 ( .I(v), .ZN(n324) );
  or2 U359 ( .A1(n325), .A2(n324), .Z(n386) );
  inv1 U361 ( .I(n353), .ZN(n326) );
  or2 U366 ( .A1(n228), .A2(n333), .Z(n401) );
  and2 U368 ( .A1(n428), .A2(n339), .Z(n340) );
  or2 U371 ( .A1(n390), .A2(g0), .Z(n345) );
  or2 U373 ( .A1(n372), .A2(q), .Z(n348) );
  and2 U374 ( .A1(n219), .A2(n350), .Z(n351) );
  or2 U376 ( .A1(n354), .A2(y), .Z(n359) );
  and2 U377 ( .A1(n428), .A2(n355), .Z(n357) );
  or2 U378 ( .A1(n249), .A2(n356), .Z(n368) );
  inv1 U381 ( .I(u), .ZN(n361) );
  and2 U383 ( .A1(s), .A2(l0), .Z(n364) );
  or2 U384 ( .A1(n364), .A2(n363), .Z(n365) );
  inv1 U385 ( .I(m), .ZN(n366) );
  or2 U386 ( .A1(n274), .A2(n366), .Z(n367) );
  and2 U387 ( .A1(k), .A2(l0), .Z(n369) );
  or2 U388 ( .A1(n369), .A2(n368), .Z(n370) );
  and2 U389 ( .A1(o), .A2(l0), .Z(n371) );
  or2 U390 ( .A1(n372), .A2(n371), .Z(n374) );
  or2 U392 ( .A1(n374), .A2(n373), .Z(n414) );
  inv1 U393 ( .I(n414), .ZN(n422) );
  or2 U395 ( .A1(n260), .A2(n375), .Z(n411) );
  inv1 U396 ( .I(n376), .ZN(n380) );
  inv1 U397 ( .I(n428), .ZN(n378) );
  inv1 U398 ( .I(i0), .ZN(n377) );
  or2 U399 ( .A1(n378), .A2(n377), .Z(n379) );
  and2 U400 ( .A1(n380), .A2(n379), .Z(n383) );
  inv1 U401 ( .I(j0), .ZN(n381) );
  inv1 U404 ( .I(y), .ZN(n384) );
  and2 U406 ( .A1(w), .A2(l0), .Z(n387) );
  or2 U407 ( .A1(n387), .A2(n386), .Z(n388) );
  or2 U408 ( .A1(n389), .A2(n262), .Z(n398) );
  and2 U409 ( .A1(e0), .A2(l0), .Z(n391) );
  or2 U410 ( .A1(n391), .A2(n390), .Z(n392) );
  or2 U411 ( .A1(n267), .A2(n392), .Z(n393) );
  and2 U413 ( .A1(a0), .A2(l0), .Z(n395) );
  or2 U414 ( .A1(n395), .A2(n394), .Z(n396) );
  or2 U417 ( .A1(n413), .A2(n420), .Z(n397) );
  inv1 U419 ( .I(i), .ZN(n399) );
  or2 U420 ( .A1(n273), .A2(n399), .Z(n400) );
  and2 U421 ( .A1(g), .A2(l0), .Z(n402) );
  or2 U422 ( .A1(n402), .A2(n401), .Z(n403) );
  and2 U425 ( .A1(c), .A2(l0), .Z(n407) );
  or2 U426 ( .A1(n407), .A2(n406), .Z(n408) );
  or2 U427 ( .A1(n229), .A2(n408), .Z(n409) );
  and2 U428 ( .A1(n410), .A2(n409), .Z(n0) );
  and2 U432 ( .A1(n414), .A2(n413), .Z(n415) );
  and2 U433 ( .A1(n416), .A2(n415), .Z(n418) );
  or2 U436 ( .A1(n427), .A2(n419), .Z(p0) );
  and2 U437 ( .A1(n420), .A2(n421), .Z(n423) );
  or2 U438 ( .A1(n423), .A2(n422), .Z(n424) );
  inv1 U212 ( .I(n273), .ZN(m0) );
  inv1f U213 ( .I(n431), .ZN(n273) );
  and2 U214 ( .A1(n219), .A2(n335), .Z(n336) );
  and2 U216 ( .A1(n219), .A2(n332), .Z(n334) );
  and2f U218 ( .A1(n367), .A2(n277), .Z(n276) );
  or2 U223 ( .A1(n319), .A2(n318), .Z(n390) );
  or2 U227 ( .A1(n336), .A2(n247), .Z(n337) );
  or2f U229 ( .A1(n427), .A2(n224), .Z(n254) );
  inv1 U230 ( .I(n412), .ZN(n427) );
  and2 U234 ( .A1(n227), .A2(n246), .Z(n226) );
  or2 U238 ( .A1(n252), .A2(n388), .Z(n251) );
  or2 U239 ( .A1(n220), .A2(n304), .Z(n347) );
  and2 U242 ( .A1(k0), .A2(f0), .Z(n323) );
  and2 U250 ( .A1(n219), .A2(n341), .Z(n342) );
  or2 U252 ( .A1(n357), .A2(n245), .Z(n358) );
  inv1 U253 ( .I(n352), .ZN(n257) );
  and2 U258 ( .A1(n385), .A2(n263), .Z(n262) );
  inv1 U261 ( .I(n393), .ZN(n420) );
  or2 U263 ( .A1(n273), .A2(n361), .Z(n362) );
  or2 U266 ( .A1(n250), .A2(n268), .Z(n207) );
  and2 U270 ( .A1(n425), .A2(n424), .Z(n426) );
  or2 U272 ( .A1(n224), .A2(n411), .Z(o0) );
  or2f U273 ( .A1(n418), .A2(n417), .Z(n419) );
  and2 U274 ( .A1(n362), .A2(n261), .Z(n260) );
  or2 U277 ( .A1(n213), .A2(n325), .Z(n353) );
  inv1 U280 ( .I(n421), .ZN(n413) );
  or2f U282 ( .A1(n292), .A2(n291), .Z(n298) );
  or2f U283 ( .A1(n342), .A2(n258), .Z(n343) );
  inv1 U285 ( .I(n343), .ZN(n269) );
  or2 U286 ( .A1(n224), .A2(n276), .Z(n417) );
  or2f U287 ( .A1(n254), .A2(n426), .Z(q0) );
  or2f U289 ( .A1(n305), .A2(n239), .Z(n315) );
  or2f U290 ( .A1(n240), .A2(n386), .Z(n354) );
  or2f U291 ( .A1(n313), .A2(n312), .Z(n314) );
  and2f U292 ( .A1(n382), .A2(n383), .Z(n389) );
  or2f U294 ( .A1(n273), .A2(n381), .Z(n382) );
  or2f U305 ( .A1(n329), .A2(n328), .Z(n330) );
  or2f U308 ( .A1(n326), .A2(n327), .Z(n328) );
  inv1f U309 ( .I(n214), .ZN(k0) );
  or2f U314 ( .A1(n260), .A2(n251), .Z(n265) );
  or2f U319 ( .A1(n242), .A2(n257), .Z(n256) );
  or2f U320 ( .A1(n271), .A2(n239), .Z(n238) );
  or2f U328 ( .A1(n405), .A2(n411), .Z(n410) );
  and2f U329 ( .A1(n431), .A2(c0), .Z(n264) );
  and2f U331 ( .A1(n431), .A2(q), .Z(n373) );
  or2f U341 ( .A1(n317), .A2(n233), .Z(n335) );
  or2f U342 ( .A1(n346), .A2(n345), .Z(n349) );
  and2f U347 ( .A1(n219), .A2(n344), .Z(n346) );
  or2f U349 ( .A1(n375), .A2(n265), .Z(n412) );
  or2f U353 ( .A1(n307), .A2(k), .Z(n355) );
  and2f U360 ( .A1(n210), .A2(n211), .Z(n307) );
  or2f U362 ( .A1(n360), .A2(n270), .Z(n231) );
  or2f U363 ( .A1(n286), .A2(n285), .Z(n287) );
  or2f U364 ( .A1(n284), .A2(n283), .Z(n286) );
  or2f U365 ( .A1(n276), .A2(n422), .Z(n375) );
  or2f U367 ( .A1(n331), .A2(n330), .Z(n219) );
  or2f U369 ( .A1(n404), .A2(n224), .Z(n405) );
  or2f U370 ( .A1(n397), .A2(n398), .Z(n404) );
  and2f U372 ( .A1(n428), .A2(n353), .Z(n240) );
  or2f U375 ( .A1(n331), .A2(n330), .Z(n428) );
  or2f U379 ( .A1(n314), .A2(n315), .Z(n331) );
  or2f U380 ( .A1(n264), .A2(n396), .Z(n421) );
  and2f U382 ( .A1(n231), .A2(g0), .Z(n267) );
  or2f U391 ( .A1(n226), .A2(n269), .Z(n268) );
  or2f U394 ( .A1(n298), .A2(n297), .Z(n299) );
  or2f U402 ( .A1(n296), .A2(n295), .Z(n297) );
  or2f U403 ( .A1(n274), .A2(n384), .Z(n385) );
  and2f U405 ( .A1(n338), .A2(n337), .Z(n248) );
  inv1f U412 ( .I(n231), .ZN(n274) );
  inv1f U415 ( .I(n219), .ZN(n271) );
  or2f U416 ( .A1(n300), .A2(n299), .Z(n222) );
  or2f U418 ( .A1(n287), .A2(n288), .Z(n300) );
  or2f U423 ( .A1(n360), .A2(n207), .Z(n431) );
  and2f U424 ( .A1(n222), .A2(b0), .Z(n319) );
  or2f U429 ( .A1(n256), .A2(n216), .Z(n360) );
endmodule

