
module i4 ( V192, V189, V186, V183, V180, V168, V156, V144, V126, V132, V88, 
        V120, V28, V56, V198, V194 );
  input [2:0] V192;
  input [2:0] V189;
  input [2:0] V186;
  input [2:0] V183;
  input [14:0] V180;
  input [14:0] V168;
  input [14:0] V156;
  input [14:0] V144;
  input [5:0] V126;
  input [5:0] V132;
  input [31:0] V88;
  input [31:0] V120;
  input [27:0] V28;
  input [27:0] V56;
  output [3:0] V198;
  output [1:0] V194;
  wire   V180_10, V180_9, V180_8, V180_6, V180_5, V180_4, V180_2, V180_1,
         V180_0, V168_10, V168_9, V168_8, V168_6, V168_5, V168_4, V168_2,
         V168_1, V168_0, V156_10, V156_9, V156_8, V156_6, V156_5, V156_4,
         V156_2, V156_1, V156_0, V144_10, V144_9, V144_8, V144_6, V144_5,
         V144_4, V144_2, V144_1, V144_0, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n40, n41, n42, n43, n44, n45, n71, n72, n73,
         n74, n75, n76, n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89,
         n90, n117, n119, n120, n121, n123, n124, n125, n126, n127, n128, n130,
         n131, n132, n133, n134, n135, n161, n162, n163, n164, n165, n166,
         n168, n169, n170, n171, n172, n173, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n198, n199, n201, n202, n205,
         n207, n208, n209, n210, n211, n212, n213, n214, n216, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n234, n235, n236, n237, n238, n240, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n259, n261, n262, n263, n264, n265, n266, n267, n268, n270, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n286, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318;
  assign V180_10 = V180[10];
  assign V180_9 = V180[9];
  assign V180_8 = V180[8];
  assign V180_6 = V180[6];
  assign V180_5 = V180[5];
  assign V180_4 = V180[4];
  assign V180_2 = V180[2];
  assign V180_1 = V180[1];
  assign V180_0 = V180[0];
  assign V168_10 = V168[10];
  assign V168_9 = V168[9];
  assign V168_8 = V168[8];
  assign V168_6 = V168[6];
  assign V168_5 = V168[5];
  assign V168_4 = V168[4];
  assign V168_2 = V168[2];
  assign V168_1 = V168[1];
  assign V168_0 = V168[0];
  assign V156_10 = V156[10];
  assign V156_9 = V156[9];
  assign V156_8 = V156[8];
  assign V156_6 = V156[6];
  assign V156_5 = V156[5];
  assign V156_4 = V156[4];
  assign V156_2 = V156[2];
  assign V156_1 = V156[1];
  assign V156_0 = V156[0];
  assign V144_10 = V144[10];
  assign V144_9 = V144[9];
  assign V144_8 = V144[8];
  assign V144_6 = V144[6];
  assign V144_5 = V144[5];
  assign V144_4 = V144[4];
  assign V144_2 = V144[2];
  assign V144_1 = V144[1];
  assign V144_0 = V144[0];

  and2f U23 ( .A1(V180_9), .A2(n28), .Z(n26) );
  and2f U26 ( .A1(n31), .A2(V180_10), .Z(n29) );
  and2f U27 ( .A1(V132[1]), .A2(V126[1]), .Z(n31) );
  and2f U69 ( .A1(V168_9), .A2(n73), .Z(n71) );
  and2f U72 ( .A1(n76), .A2(V88[17]), .Z(n74) );
  and2f U73 ( .A1(V168_10), .A2(V120[17]), .Z(n76) );
  and2f U114 ( .A1(V56[27]), .A2(V28[27]), .Z(n117) );
  and2f U117 ( .A1(V88[0]), .A2(V120[0]), .Z(n120) );
  and2f U118 ( .A1(n121), .A2(V88[1]), .Z(n119) );
  and2f U119 ( .A1(V156_10), .A2(V120[1]), .Z(n121) );
  and2f U127 ( .A1(n128), .A2(V56[25]), .Z(n126) );
  and2f U128 ( .A1(V28[25]), .A2(V156_6), .Z(n128) );
  and2f U161 ( .A1(V144_9), .A2(n163), .Z(n161) );
  and2f U164 ( .A1(n166), .A2(V56[13]), .Z(n164) );
  and2f U165 ( .A1(V28[13]), .A2(V144_10), .Z(n166) );
  and2f U170 ( .A1(V144_5), .A2(n170), .Z(n168) );
  and2f U173 ( .A1(n173), .A2(V56[9]), .Z(n171) );
  and2f U174 ( .A1(V28[9]), .A2(V144_6), .Z(n173) );
  and2f U191 ( .A1(V28[17]), .A2(V144[14]), .Z(n182) );
  and2f U192 ( .A1(n182), .A2(V56[17]), .Z(n184) );
  or2f U194 ( .A1(n184), .A2(n183), .Z(n185) );
  and2f U195 ( .A1(n185), .A2(V144[13]), .Z(n187) );
  or2f U197 ( .A1(n187), .A2(n186), .Z(n188) );
  and2f U198 ( .A1(n188), .A2(V144[12]), .Z(n190) );
  or2f U200 ( .A1(n190), .A2(n189), .Z(n191) );
  and2f U201 ( .A1(n191), .A2(V183[2]), .Z(n196) );
  or2f U202 ( .A1(n161), .A2(n162), .Z(n192) );
  and2f U203 ( .A1(n192), .A2(V144_8), .Z(n194) );
  and2f U219 ( .A1(V88[5]), .A2(V156[14]), .Z(n209) );
  and2f U220 ( .A1(n209), .A2(V120[5]), .Z(n211) );
  or2f U222 ( .A1(n211), .A2(n210), .Z(n212) );
  and2f U223 ( .A1(n212), .A2(V156[13]), .Z(n214) );
  and2f U231 ( .A1(n219), .A2(V156_8), .Z(n221) );
  or2f U233 ( .A1(n221), .A2(n220), .Z(n222) );
  or2f U234 ( .A1(n223), .A2(n222), .Z(n224) );
  and2f U235 ( .A1(n224), .A2(V186[1]), .Z(n227) );
  or2f U238 ( .A1(n227), .A2(n226), .Z(n228) );
  or2f U239 ( .A1(n229), .A2(n228), .Z(n230) );
  and2f U240 ( .A1(n230), .A2(V186[0]), .Z(n231) );
  or2f U242 ( .A1(n231), .A2(n303), .Z(V198[1]) );
  and2f U247 ( .A1(V88[21]), .A2(V168[14]), .Z(n236) );
  and2f U248 ( .A1(n236), .A2(V120[21]), .Z(n238) );
  and2f U249 ( .A1(V120[20]), .A2(V88[20]), .Z(n237) );
  and2f U252 ( .A1(V120[19]), .A2(V88[19]), .Z(n240) );
  and2f U254 ( .A1(n242), .A2(V168[12]), .Z(n244) );
  or2f U256 ( .A1(n244), .A2(n243), .Z(n245) );
  and2f U257 ( .A1(n245), .A2(V189[2]), .Z(n250) );
  or2f U258 ( .A1(n71), .A2(n72), .Z(n246) );
  and2f U259 ( .A1(n246), .A2(V168_8), .Z(n248) );
  or2f U262 ( .A1(n250), .A2(n249), .Z(n251) );
  and2f U263 ( .A1(n251), .A2(V189[1]), .Z(n254) );
  or2f U266 ( .A1(n254), .A2(n253), .Z(n255) );
  and2f U275 ( .A1(V126[5]), .A2(V180[14]), .Z(n263) );
  and2f U276 ( .A1(n263), .A2(V132[5]), .Z(n265) );
  or2f U278 ( .A1(n265), .A2(n264), .Z(n266) );
  and2f U279 ( .A1(n266), .A2(V180[13]), .Z(n268) );
  and2f U285 ( .A1(n272), .A2(V192[2]), .Z(n277) );
  or2f U286 ( .A1(n26), .A2(n27), .Z(n273) );
  and2f U287 ( .A1(n273), .A2(V180_8), .Z(n275) );
  or2f U290 ( .A1(n277), .A2(n276), .Z(n278) );
  and2f U291 ( .A1(n278), .A2(V192[1]), .Z(n281) );
  or2f U294 ( .A1(n281), .A2(n280), .Z(n282) );
  and2 U187 ( .A1(V56[11]), .A2(V28[11]), .Z(n162) );
  and2 U188 ( .A1(V88[15]), .A2(V120[15]), .Z(n72) );
  and2 U189 ( .A1(V88[31]), .A2(V120[31]), .Z(n27) );
  or2f U190 ( .A1(n194), .A2(n193), .Z(n195) );
  or2f U193 ( .A1(n248), .A2(n247), .Z(n249) );
  or2f U196 ( .A1(n275), .A2(n274), .Z(n276) );
  and2 U199 ( .A1(V120[4]), .A2(V88[4]), .Z(n210) );
  and2 U204 ( .A1(V180_6), .A2(V120[29]), .Z(n38) );
  or2 U205 ( .A1(n267), .A2(n270), .Z(n318) );
  and2 U206 ( .A1(n83), .A2(V88[13]), .Z(n81) );
  and2 U207 ( .A1(V168_6), .A2(V120[13]), .Z(n83) );
  and2 U208 ( .A1(V132[3]), .A2(V126[3]), .Z(n267) );
  and2 U209 ( .A1(V132[4]), .A2(V126[4]), .Z(n264) );
  or2 U210 ( .A1(n29), .A2(n30), .Z(n28) );
  and2 U211 ( .A1(V132[0]), .A2(V126[0]), .Z(n30) );
  or2 U212 ( .A1(n164), .A2(n165), .Z(n163) );
  and2 U213 ( .A1(V56[12]), .A2(V28[12]), .Z(n165) );
  and2 U214 ( .A1(V56[16]), .A2(V28[16]), .Z(n183) );
  and2 U215 ( .A1(V56[15]), .A2(V28[15]), .Z(n186) );
  or2 U216 ( .A1(n213), .A2(n216), .Z(n311) );
  and2 U217 ( .A1(V120[3]), .A2(V88[3]), .Z(n213) );
  or2 U218 ( .A1(n74), .A2(n75), .Z(n73) );
  and2 U221 ( .A1(V88[16]), .A2(V120[16]), .Z(n75) );
  and2 U224 ( .A1(V156_5), .A2(n125), .Z(n123) );
  and2 U225 ( .A1(V180_5), .A2(n35), .Z(n33) );
  and2 U226 ( .A1(n38), .A2(V88[29]), .Z(n36) );
  and2 U227 ( .A1(V168_5), .A2(n80), .Z(n78) );
  or2f U228 ( .A1(n119), .A2(n291), .Z(n289) );
  and2f U229 ( .A1(n289), .A2(n290), .Z(n219) );
  or2 U230 ( .A1(n117), .A2(V156_9), .Z(n290) );
  or2f U232 ( .A1(n120), .A2(n117), .Z(n291) );
  or2f U236 ( .A1(n196), .A2(n294), .Z(n292) );
  and2f U237 ( .A1(n292), .A2(n293), .Z(n201) );
  or2 U241 ( .A1(n199), .A2(V183[1]), .Z(n293) );
  or2f U243 ( .A1(n195), .A2(n199), .Z(n294) );
  and2f U244 ( .A1(n198), .A2(V144_4), .Z(n199) );
  or2f U245 ( .A1(n238), .A2(n297), .Z(n295) );
  and2f U246 ( .A1(n295), .A2(n296), .Z(n242) );
  or2 U250 ( .A1(n240), .A2(V168[13]), .Z(n296) );
  or2f U251 ( .A1(n237), .A2(n240), .Z(n297) );
  or2 U253 ( .A1(n214), .A2(n311), .Z(n298) );
  and2f U255 ( .A1(n298), .A2(n299), .Z(n223) );
  and2 U260 ( .A1(V186[2]), .A2(n310), .Z(n299) );
  or2f U261 ( .A1(n282), .A2(n302), .Z(n300) );
  and2f U264 ( .A1(n300), .A2(n301), .Z(V198[3]) );
  or2 U265 ( .A1(n288), .A2(n304), .Z(n301) );
  or2f U267 ( .A1(n305), .A2(n288), .Z(n302) );
  and2f U268 ( .A1(V144_0), .A2(n181), .Z(n205) );
  or2f U269 ( .A1(n175), .A2(n176), .Z(n181) );
  and2f U270 ( .A1(V168_0), .A2(n235), .Z(n259) );
  or2f U271 ( .A1(n85), .A2(n86), .Z(n235) );
  and2f U272 ( .A1(n45), .A2(V88[25]), .Z(n43) );
  and2f U273 ( .A1(V180_0), .A2(n262), .Z(n286) );
  or2 U274 ( .A1(n232), .A2(n234), .Z(n303) );
  or2 U277 ( .A1(n286), .A2(V192[0]), .Z(n304) );
  or2f U280 ( .A1(n283), .A2(n286), .Z(n305) );
  or2f U281 ( .A1(n205), .A2(n207), .Z(n306) );
  or2f U282 ( .A1(n201), .A2(n309), .Z(n307) );
  and2f U283 ( .A1(n307), .A2(n308), .Z(V198[0]) );
  or2 U284 ( .A1(n306), .A2(V183[0]), .Z(n308) );
  or2f U288 ( .A1(n202), .A2(n306), .Z(n309) );
  or2 U289 ( .A1(n216), .A2(V156[12]), .Z(n310) );
  or2f U292 ( .A1(n259), .A2(n261), .Z(n312) );
  or2f U293 ( .A1(n255), .A2(n315), .Z(n313) );
  and2f U295 ( .A1(n313), .A2(n314), .Z(V198[2]) );
  or2 U296 ( .A1(n312), .A2(V189[0]), .Z(n314) );
  or2f U297 ( .A1(n256), .A2(n312), .Z(n315) );
  or2f U298 ( .A1(n268), .A2(n318), .Z(n316) );
  and2f U299 ( .A1(n316), .A2(n317), .Z(n272) );
  or2 U300 ( .A1(n270), .A2(V180[12]), .Z(n317) );
  or2 U301 ( .A1(n171), .A2(n172), .Z(n170) );
  and2 U302 ( .A1(V56[8]), .A2(V28[8]), .Z(n172) );
  or2 U303 ( .A1(n126), .A2(n127), .Z(n125) );
  and2 U304 ( .A1(V56[24]), .A2(V28[24]), .Z(n127) );
  or2 U305 ( .A1(n81), .A2(n82), .Z(n80) );
  and2 U306 ( .A1(V88[12]), .A2(V120[12]), .Z(n82) );
  or2 U307 ( .A1(n36), .A2(n37), .Z(n35) );
  and2 U308 ( .A1(V88[28]), .A2(V120[28]), .Z(n37) );
  and2 U309 ( .A1(V56[3]), .A2(V28[3]), .Z(n176) );
  and2 U310 ( .A1(V144_1), .A2(n177), .Z(n175) );
  or2 U311 ( .A1(n178), .A2(n179), .Z(n177) );
  and2 U312 ( .A1(V56[6]), .A2(V28[6]), .Z(n202) );
  or2 U313 ( .A1(n130), .A2(n131), .Z(n208) );
  and2 U314 ( .A1(V56[19]), .A2(V28[19]), .Z(n131) );
  and2 U315 ( .A1(V156_1), .A2(n132), .Z(n130) );
  or2 U316 ( .A1(n133), .A2(n134), .Z(n132) );
  and2 U317 ( .A1(V56[22]), .A2(V28[22]), .Z(n229) );
  and2 U318 ( .A1(V88[7]), .A2(V120[7]), .Z(n86) );
  and2 U319 ( .A1(V168_1), .A2(n87), .Z(n85) );
  or2 U320 ( .A1(n88), .A2(n89), .Z(n87) );
  and2 U321 ( .A1(V120[10]), .A2(V88[10]), .Z(n256) );
  or2 U322 ( .A1(n40), .A2(n41), .Z(n262) );
  and2 U323 ( .A1(V88[23]), .A2(V120[23]), .Z(n41) );
  and2 U324 ( .A1(V180_1), .A2(n42), .Z(n40) );
  or2 U325 ( .A1(n43), .A2(n44), .Z(n42) );
  and2 U326 ( .A1(V120[26]), .A2(V88[26]), .Z(n283) );
  and2 U327 ( .A1(V56[14]), .A2(V28[14]), .Z(n189) );
  and2 U328 ( .A1(V56[10]), .A2(V28[10]), .Z(n193) );
  and2 U329 ( .A1(V120[2]), .A2(V88[2]), .Z(n216) );
  and2 U330 ( .A1(V56[26]), .A2(V28[26]), .Z(n220) );
  and2 U331 ( .A1(V120[18]), .A2(V88[18]), .Z(n243) );
  and2 U332 ( .A1(V120[14]), .A2(V88[14]), .Z(n247) );
  and2 U333 ( .A1(V132[2]), .A2(V126[2]), .Z(n270) );
  and2 U334 ( .A1(V120[30]), .A2(V88[30]), .Z(n274) );
  and2 U335 ( .A1(n180), .A2(V56[5]), .Z(n178) );
  and2 U336 ( .A1(V28[5]), .A2(V144_2), .Z(n180) );
  and2 U337 ( .A1(V56[4]), .A2(V28[4]), .Z(n179) );
  or2 U338 ( .A1(n168), .A2(n169), .Z(n198) );
  and2 U339 ( .A1(V56[7]), .A2(V28[7]), .Z(n169) );
  and2 U340 ( .A1(n135), .A2(V56[21]), .Z(n133) );
  and2 U341 ( .A1(V28[21]), .A2(V156_2), .Z(n135) );
  and2 U342 ( .A1(V56[20]), .A2(V28[20]), .Z(n134) );
  and2 U343 ( .A1(n225), .A2(V156_4), .Z(n226) );
  or2 U344 ( .A1(n123), .A2(n124), .Z(n225) );
  and2 U345 ( .A1(V56[23]), .A2(V28[23]), .Z(n124) );
  and2 U346 ( .A1(n90), .A2(V88[9]), .Z(n88) );
  and2 U347 ( .A1(V168_2), .A2(V120[9]), .Z(n90) );
  and2 U348 ( .A1(V88[8]), .A2(V120[8]), .Z(n89) );
  and2 U349 ( .A1(n252), .A2(V168_4), .Z(n253) );
  or2 U350 ( .A1(n78), .A2(n79), .Z(n252) );
  and2 U351 ( .A1(V88[11]), .A2(V120[11]), .Z(n79) );
  and2 U352 ( .A1(V180_2), .A2(V120[25]), .Z(n45) );
  and2 U353 ( .A1(V88[24]), .A2(V120[24]), .Z(n44) );
  and2 U354 ( .A1(n279), .A2(V180_4), .Z(n280) );
  or2 U355 ( .A1(n33), .A2(n34), .Z(n279) );
  and2 U356 ( .A1(V88[27]), .A2(V120[27]), .Z(n34) );
  and2 U357 ( .A1(V28[2]), .A2(V56[2]), .Z(n207) );
  and2 U358 ( .A1(V28[18]), .A2(V56[18]), .Z(n234) );
  and2 U359 ( .A1(V156_0), .A2(n208), .Z(n232) );
  and2 U360 ( .A1(V88[6]), .A2(V120[6]), .Z(n261) );
  and2 U361 ( .A1(V88[22]), .A2(V120[22]), .Z(n288) );
  and2 U362 ( .A1(V56[0]), .A2(V28[0]), .Z(V194[0]) );
  and2 U363 ( .A1(V56[1]), .A2(V28[1]), .Z(V194[1]) );
endmodule

