
module pair ( r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, 
        b5, a5, z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, 
        j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, 
        r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, 
        z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2, 
        h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1, 
        p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0, y0, 
        x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0, h0, g0, 
        f0, e0, d0, c0, b0, a0, z, y, w, v, u, t, s, r, q, p, o, n, m, l, k, j, 
        i, h, g, f, e, d, c, b, a, y10, x10, w10, v10, u10, t10, s10, r10, q10, 
        p10, o10, n10, m10, l10, k10, j10, i10, h10, g10, f10, e10, d10, c10, 
        b10, a10, z9, y9, x9, w9, v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, 
        k9, j9, i9, h9, g9, f9, e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8, 
        s8, r8, q8, p8, o8, n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8, b8, 
        a8, z7, y7, x7, w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, 
        i7, h7, g7, f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, 
        q6, p6, o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, 
        y5, x5, w5, v5, u5, t5, s5 );
  input r5, q5, p5, o5, n5, m5, l5, k5, j5, i5, h5, g5, f5, e5, d5, c5, b5, a5,
         z4, y4, x4, w4, v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4,
         i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3,
         r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3,
         a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2,
         j2, i2, h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1,
         s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1,
         b1, a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0,
         k0, j0, i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, w, v, u, t, s, r, q,
         p, o, n, m, l, k, j, i, h, g, f, e, d, c, b, a;
  output y10, x10, w10, v10, u10, t10, s10, r10, q10, p10, o10, n10, m10, l10,
         k10, j10, i10, h10, g10, f10, e10, d10, c10, b10, a10, z9, y9, x9, w9,
         v9, u9, t9, s9, r9, q9, p9, o9, n9, m9, l9, k9, j9, i9, h9, g9, f9,
         e9, d9, c9, b9, a9, z8, y8, x8, w8, v8, u8, t8, s8, r8, q8, p8, o8,
         n8, m8, l8, k8, j8, i8, h8, g8, f8, e8, d8, c8, b8, a8, z7, y7, x7,
         w7, v7, u7, t7, s7, r7, q7, p7, o7, n7, m7, l7, k7, j7, i7, h7, g7,
         f7, e7, d7, c7, b7, a7, z6, y6, x6, w6, v6, u6, t6, s6, r6, q6, p6,
         o6, n6, m6, l6, k6, j6, i6, h6, g6, f6, e6, d6, c6, b6, a6, z5, y5,
         x5, w5, v5, u5, t5, s5;
  wire   n1966, n1967, n1968, n1969, n1970, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n323, n324, n325, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n653, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n742, n743, n745, n746, n747, n748, n749, n750, n751, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n915, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n952, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1047, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1060, n1061, n1062, n1063, n1065, n1068, n1070,
         n1071, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1089, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1203,
         n1205, n1206, n1207, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1258, n1261, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1447,
         n1454, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1481, n1482, n1483, n1484, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1548, n1549, n1550, n1551, n1552, n1554, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1603, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1617, n1618, n1619, n1620,
         n1621, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1690, n1692, n1696, n1698, n1699,
         n1715, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1742, n1743, n1744, n1745, n1746,
         n1747, n1749, n1750, n1751, n1754, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1894, n1895, n1896, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1945,
         n1946, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068;

  or2f U5 ( .A1(n245), .A2(n246), .Z(z8) );
  and2f U6 ( .A1(n247), .A2(n248), .Z(n245) );
  or2f U7 ( .A1(n249), .A2(n250), .Z(n248) );
  and2f U8 ( .A1(n251), .A2(n252), .Z(n250) );
  inv1f U9 ( .I(n253), .ZN(n251) );
  or2f U11 ( .A1(n255), .A2(n254), .Z(n253) );
  or2f U12 ( .A1(n256), .A2(n257), .Z(n255) );
  and2f U14 ( .A1(n259), .A2(n260), .Z(n256) );
  and2f U15 ( .A1(n261), .A2(n262), .Z(z7) );
  or2f U16 ( .A1(n263), .A2(n264), .Z(n262) );
  or2f U18 ( .A1(n266), .A2(s2), .Z(n265) );
  and2f U19 ( .A1(s2), .A2(n266), .Z(n263) );
  or2f U20 ( .A1(n267), .A2(n268), .Z(n266) );
  and2f U57 ( .A1(n312), .A2(n313), .Z(n311) );
  or2f U58 ( .A1(n314), .A2(n315), .Z(n313) );
  or2f U59 ( .A1(r3), .A2(n316), .Z(n315) );
  and2f U60 ( .A1(n317), .A2(n318), .Z(n316) );
  and2f U68 ( .A1(n328), .A2(n329), .Z(n327) );
  and2f U71 ( .A1(r2), .A2(n330), .Z(n331) );
  or2f U73 ( .A1(n334), .A2(n335), .Z(n332) );
  and2f U74 ( .A1(n2023), .A2(n336), .Z(n335) );
  or2f U115 ( .A1(n383), .A2(z), .Z(x9) );
  and2f U116 ( .A1(n384), .A2(n385), .Z(n383) );
  or2f U117 ( .A1(n386), .A2(n387), .Z(n385) );
  or2f U118 ( .A1(n388), .A2(n389), .Z(n387) );
  and2f U121 ( .A1(q4), .A2(n391), .Z(n388) );
  or2f U122 ( .A1(n392), .A2(n393), .Z(n391) );
  and2f U125 ( .A1(n247), .A2(n396), .Z(n395) );
  or2f U126 ( .A1(n397), .A2(n398), .Z(n396) );
  and2f U127 ( .A1(q3), .A2(n399), .Z(n398) );
  or2f U128 ( .A1(n400), .A2(n401), .Z(n399) );
  or2f U191 ( .A1(n460), .A2(n246), .Z(w8) );
  and2f U192 ( .A1(n247), .A2(n461), .Z(n460) );
  or2f U193 ( .A1(n462), .A2(n463), .Z(n461) );
  or2f U195 ( .A1(n465), .A2(p3), .Z(n464) );
  or2f U197 ( .A1(n466), .A2(n467), .Z(n465) );
  and2f U200 ( .A1(n471), .A2(n472), .Z(n468) );
  or2f U240 ( .A1(n510), .A2(n511), .Z(n509) );
  or2f U241 ( .A1(n512), .A2(n513), .Z(n511) );
  or2f U273 ( .A1(n386), .A2(n542), .Z(n541) );
  or2f U274 ( .A1(n543), .A2(n544), .Z(n542) );
  inv1f U278 ( .I(n545), .ZN(n393) );
  and2f U279 ( .A1(n4), .A2(n546), .Z(n545) );
  and2f U286 ( .A1(o3), .A2(n552), .Z(n549) );
  or2f U287 ( .A1(n553), .A2(n554), .Z(n552) );
  or2f U288 ( .A1(n1972), .A2(n555), .Z(n554) );
  or2f U290 ( .A1(n557), .A2(n558), .Z(n556) );
  or2f U294 ( .A1(n563), .A2(b), .Z(v7) );
  and2f U295 ( .A1(n564), .A2(n565), .Z(n563) );
  or2f U296 ( .A1(n566), .A2(n567), .Z(n565) );
  or2f U297 ( .A1(n568), .A2(n569), .Z(n567) );
  inv1f U298 ( .I(n570), .ZN(n569) );
  or2f U299 ( .A1(n571), .A2(o2), .Z(n570) );
  and2f U300 ( .A1(o2), .A2(n571), .Z(n568) );
  or2f U301 ( .A1(n572), .A2(n573), .Z(n571) );
  and2f U334 ( .A1(n606), .A2(n557), .Z(n605) );
  inv1f U335 ( .I(n607), .ZN(n606) );
  or2f U337 ( .A1(n466), .A2(n608), .Z(n607) );
  and2f U385 ( .A1(n661), .A2(m4), .Z(n546) );
  or2f U387 ( .A1(n662), .A2(j0), .Z(n661) );
  and2f U388 ( .A1(n663), .A2(l4), .Z(n662) );
  and2f U389 ( .A1(n664), .A2(k4), .Z(n663) );
  and2f U392 ( .A1(n666), .A2(n667), .Z(n665) );
  or2f U393 ( .A1(n668), .A2(n669), .Z(n667) );
  or2f U394 ( .A1(m3), .A2(n670), .Z(n669) );
  and2f U395 ( .A1(n671), .A2(n672), .Z(n670) );
  and2f U396 ( .A1(n2049), .A2(n673), .Z(n671) );
  or2f U408 ( .A1(n566), .A2(n682), .Z(n681) );
  or2f U409 ( .A1(n683), .A2(n684), .Z(n682) );
  inv1f U413 ( .I(n685), .ZN(n572) );
  and2f U414 ( .A1(n2020), .A2(n836), .Z(n685) );
  and2f U494 ( .A1(n772), .A2(n773), .Z(n771) );
  or2f U495 ( .A1(n774), .A2(n775), .Z(n773) );
  or2f U496 ( .A1(l3), .A2(n776), .Z(n775) );
  or2f U504 ( .A1(n780), .A2(n402), .Z(n466) );
  or2f U509 ( .A1(n781), .A2(b), .Z(s7) );
  or2f U511 ( .A1(n566), .A2(n784), .Z(n783) );
  and2f U560 ( .A1(h4), .A2(n826), .Z(n664) );
  and2f U561 ( .A1(j4), .A2(n827), .Z(n826) );
  and2f U572 ( .A1(n836), .A2(k2), .Z(n686) );
  or2f U574 ( .A1(n837), .A2(l), .Z(n836) );
  and2f U575 ( .A1(n838), .A2(j2), .Z(n837) );
  and2f U576 ( .A1(i2), .A2(n839), .Z(n838) );
  and2f U629 ( .A1(n247), .A2(n891), .Z(n890) );
  or2f U630 ( .A1(n892), .A2(n893), .Z(n891) );
  or2f U632 ( .A1(n895), .A2(i3), .Z(n894) );
  or2f U636 ( .A1(n899), .A2(n2037), .Z(n898) );
  and2f U647 ( .A1(h2), .A2(n908), .Z(n839) );
  and2f U648 ( .A1(n909), .A2(f2), .Z(n908) );
  or2f U665 ( .A1(n926), .A2(n927), .Z(n925) );
  or2f U667 ( .A1(n929), .A2(h3), .Z(n928) );
  or2f U669 ( .A1(n930), .A2(n931), .Z(n929) );
  or2f U706 ( .A1(n968), .A2(n969), .Z(n967) );
  and2f U744 ( .A1(n1967), .A2(n1004), .Z(n982) );
  or2f U748 ( .A1(n1007), .A2(n1008), .Z(n1006) );
  and2f U749 ( .A1(n960), .A2(n1004), .Z(n1008) );
  or2f U759 ( .A1(n1017), .A2(n1018), .Z(l8) );
  and2f U760 ( .A1(n261), .A2(n1019), .Z(n1017) );
  or2f U761 ( .A1(n1020), .A2(n1021), .Z(n1019) );
  or2f U763 ( .A1(n1023), .A2(e3), .Z(n1022) );
  or2f U765 ( .A1(n1025), .A2(n1024), .Z(n1023) );
  or2f U766 ( .A1(n1026), .A2(n1027), .Z(n1025) );
  and2f U769 ( .A1(n1028), .A2(n1978), .Z(n1026) );
  or2f U770 ( .A1(n1029), .A2(n1030), .Z(n1028) );
  and2f U781 ( .A1(n1036), .A2(e2), .Z(n909) );
  or2f U782 ( .A1(n974), .A2(n1037), .Z(n1036) );
  and2f U784 ( .A1(n975), .A2(g2), .Z(n974) );
  or2f U785 ( .A1(n1038), .A2(n1039), .Z(n975) );
  or2f U795 ( .A1(n1049), .A2(n1018), .Z(k8) );
  and2f U796 ( .A1(n261), .A2(n1050), .Z(n1049) );
  or2f U797 ( .A1(n1051), .A2(n1052), .Z(n1050) );
  and2f U798 ( .A1(n1053), .A2(n1029), .Z(n1052) );
  or2f U802 ( .A1(n1024), .A2(n1055), .Z(n1054) );
  or2f U803 ( .A1(n1056), .A2(n1057), .Z(n1055) );
  and2f U804 ( .A1(c3), .A2(n2023), .Z(n1057) );
  and2f U805 ( .A1(n1978), .A2(n1030), .Z(n1056) );
  or2f U806 ( .A1(n2046), .A2(n2042), .Z(n1030) );
  and2f U810 ( .A1(d2), .A2(n1063), .Z(n1039) );
  and2f U812 ( .A1(c2), .A2(b2), .Z(n1063) );
  or2f U824 ( .A1(n1075), .A2(n1076), .Z(j9) );
  and2f U826 ( .A1(n1078), .A2(n1079), .Z(n1077) );
  or2f U827 ( .A1(n1080), .A2(n1081), .Z(n1078) );
  or2f U829 ( .A1(n1083), .A2(c4), .Z(n1082) );
  and2f U830 ( .A1(c4), .A2(n1083), .Z(n1080) );
  or2f U831 ( .A1(n1084), .A2(n1085), .Z(n1083) );
  or2f U832 ( .A1(n1086), .A2(n1087), .Z(n1085) );
  and2f U837 ( .A1(n1094), .A2(n261), .Z(j8) );
  and2f U838 ( .A1(n1095), .A2(n1096), .Z(n1094) );
  or2f U839 ( .A1(n1097), .A2(n1098), .Z(n1096) );
  or2f U840 ( .A1(c3), .A2(n1099), .Z(n1098) );
  and2f U841 ( .A1(n1100), .A2(n1101), .Z(n1099) );
  or2f U849 ( .A1(n1107), .A2(n269), .Z(n1024) );
  and2f U850 ( .A1(n2022), .A2(n1108), .Z(n1107) );
  or2f U861 ( .A1(n1117), .A2(n1118), .Z(i9) );
  and2f U863 ( .A1(n1120), .A2(n1079), .Z(n1119) );
  or2f U864 ( .A1(n1121), .A2(n1122), .Z(n1120) );
  and2f U865 ( .A1(n1123), .A2(n1091), .Z(n1122) );
  inv1f U867 ( .I(n1124), .ZN(n1123) );
  and2f U868 ( .A1(b4), .A2(n1124), .Z(n1121) );
  or2f U869 ( .A1(n1125), .A2(n1084), .Z(n1124) );
  or2f U870 ( .A1(n1126), .A2(n1127), .Z(n1084) );
  or2f U875 ( .A1(n1130), .A2(n1018), .Z(i8) );
  and2f U876 ( .A1(n261), .A2(n1131), .Z(n1130) );
  or2f U877 ( .A1(n1132), .A2(n1133), .Z(n1131) );
  and2f U878 ( .A1(b3), .A2(n1134), .Z(n1133) );
  or2f U879 ( .A1(n1135), .A2(n1136), .Z(n1134) );
  or2f U894 ( .A1(n2022), .A2(n1106), .Z(n1138) );
  or2f U895 ( .A1(n1149), .A2(j), .Z(n1106) );
  and2f U896 ( .A1(n1150), .A2(v2), .Z(n1149) );
  or2f U914 ( .A1(n1166), .A2(n1167), .Z(n1127) );
  or2f U923 ( .A1(n1177), .A2(n1018), .Z(h8) );
  and2f U924 ( .A1(n261), .A2(n1178), .Z(n1177) );
  or2f U925 ( .A1(n1179), .A2(n1180), .Z(n1178) );
  inv1f U926 ( .I(n1181), .ZN(n1180) );
  or2f U927 ( .A1(n1182), .A2(a3), .Z(n1181) );
  and2f U928 ( .A1(a3), .A2(n1182), .Z(n1179) );
  or2f U929 ( .A1(n1183), .A2(n1184), .Z(n1182) );
  and2f U931 ( .A1(n1186), .A2(n1187), .Z(n1185) );
  or2f U933 ( .A1(n1188), .A2(n2023), .Z(n1186) );
  or2f U935 ( .A1(n1189), .A2(n1190), .Z(h7) );
  or2f U936 ( .A1(b), .A2(n1191), .Z(n1190) );
  and2f U937 ( .A1(n1192), .A2(n1193), .Z(n1191) );
  or2f U938 ( .A1(n1194), .A2(n1195), .Z(n1192) );
  or2f U940 ( .A1(n1197), .A2(a2), .Z(n1196) );
  or2f U942 ( .A1(n1198), .A2(n1199), .Z(n1197) );
  or2f U953 ( .A1(n1212), .A2(n1213), .Z(g9) );
  and2f U955 ( .A1(n1215), .A2(n1079), .Z(n1214) );
  or2f U956 ( .A1(n1216), .A2(n1217), .Z(n1215) );
  and2f U957 ( .A1(n1218), .A2(n1176), .Z(n1217) );
  or2f U961 ( .A1(n1220), .A2(n1221), .Z(n1219) );
  or2f U967 ( .A1(n1226), .A2(n1018), .Z(g8) );
  and2f U968 ( .A1(n261), .A2(n1227), .Z(n1226) );
  or2f U969 ( .A1(n1228), .A2(n1229), .Z(n1227) );
  inv1f U970 ( .I(n1230), .ZN(n1229) );
  or2f U971 ( .A1(n1231), .A2(z2), .Z(n1230) );
  or2f U973 ( .A1(n1232), .A2(n1233), .Z(n1231) );
  or2f U974 ( .A1(n269), .A2(n1234), .Z(n1233) );
  or2f U976 ( .A1(n703), .A2(n1236), .Z(n1235) );
  or2f U978 ( .A1(n1238), .A2(n1239), .Z(n1237) );
  or2f U980 ( .A1(n1240), .A2(n1241), .Z(g7) );
  or2f U981 ( .A1(b), .A2(n1242), .Z(n1241) );
  and2f U982 ( .A1(n1243), .A2(n1193), .Z(n1242) );
  or2f U983 ( .A1(n1244), .A2(n1245), .Z(n1243) );
  and2f U984 ( .A1(n1246), .A2(n1205), .Z(n1245) );
  inv1f U986 ( .I(n1247), .ZN(n1246) );
  or2f U988 ( .A1(n1248), .A2(n1198), .Z(n1247) );
  or2f U989 ( .A1(n1250), .A2(n1249), .Z(n1198) );
  or2f U1005 ( .A1(n1263), .A2(n1264), .Z(f9) );
  and2f U1007 ( .A1(n1266), .A2(n1079), .Z(n1265) );
  or2f U1008 ( .A1(n1267), .A2(n1268), .Z(n1266) );
  and2f U1009 ( .A1(n1269), .A2(n1224), .Z(n1268) );
  inv1f U1011 ( .I(n1270), .ZN(n1269) );
  and2f U1012 ( .A1(y3), .A2(n1270), .Z(n1267) );
  or2f U1013 ( .A1(n1271), .A2(n1220), .Z(n1270) );
  or2f U1014 ( .A1(n1272), .A2(n1273), .Z(n1220) );
  and2f U1021 ( .A1(n1279), .A2(n703), .Z(n1278) );
  and2f U1023 ( .A1(y2), .A2(n1280), .Z(n1277) );
  or2f U1024 ( .A1(n1183), .A2(n1281), .Z(n1280) );
  or2f U1025 ( .A1(n1282), .A2(n1283), .Z(n1281) );
  or2f U1027 ( .A1(n1284), .A2(n1285), .Z(n1236) );
  or2f U1038 ( .A1(n1294), .A2(n285), .Z(n1250) );
  or2f U1061 ( .A1(n1319), .A2(n1320), .Z(n1318) );
  and2f U1062 ( .A1(n1321), .A2(n1275), .Z(n1320) );
  or2f U1067 ( .A1(n1324), .A2(n1167), .Z(n1273) );
  and2f U1078 ( .A1(n1330), .A2(n261), .Z(e8) );
  and2f U1079 ( .A1(n1331), .A2(n1332), .Z(n1330) );
  or2f U1080 ( .A1(n1333), .A2(n1334), .Z(n1332) );
  or2f U1081 ( .A1(x2), .A2(n1335), .Z(n1334) );
  and2f U1082 ( .A1(n1336), .A2(n1100), .Z(n1335) );
  and2f U1084 ( .A1(n1339), .A2(n1102), .Z(n1333) );
  inv1f U1091 ( .I(n1339), .ZN(n1285) );
  and2f U1092 ( .A1(n1151), .A2(w2), .Z(n1339) );
  or2f U1093 ( .A1(n1344), .A2(n1345), .Z(e7) );
  or2f U1094 ( .A1(b), .A2(n1346), .Z(n1345) );
  and2f U1095 ( .A1(n1347), .A2(n1193), .Z(n1346) );
  or2f U1096 ( .A1(n1348), .A2(n1349), .Z(n1347) );
  and2f U1097 ( .A1(n1350), .A2(n1303), .Z(n1349) );
  inv1f U1099 ( .I(n1351), .ZN(n1350) );
  or2f U1101 ( .A1(n1352), .A2(n1353), .Z(n1351) );
  or2f U1122 ( .A1(n1371), .A2(w3), .Z(n1370) );
  or2f U1124 ( .A1(n1372), .A2(n1373), .Z(n1371) );
  and2f U1131 ( .A1(n1377), .A2(n261), .Z(d8) );
  and2f U1132 ( .A1(n1378), .A2(n1379), .Z(n1377) );
  or2f U1133 ( .A1(n1380), .A2(n1381), .Z(n1379) );
  or2f U1134 ( .A1(w2), .A2(n1382), .Z(n1381) );
  and2f U1135 ( .A1(n1100), .A2(n1337), .Z(n1382) );
  or2f U1145 ( .A1(n1386), .A2(j), .Z(n1151) );
  or2f U1147 ( .A1(n1388), .A2(n269), .Z(n1183) );
  and2f U1148 ( .A1(n1147), .A2(n2023), .Z(n1388) );
  or2f U1150 ( .A1(n1390), .A2(t2), .Z(n1389) );
  or2f U1152 ( .A1(b), .A2(n1393), .Z(n1392) );
  and2f U1153 ( .A1(n1394), .A2(n1193), .Z(n1393) );
  or2f U1154 ( .A1(n1395), .A2(n1396), .Z(n1394) );
  and2f U1155 ( .A1(n1397), .A2(n1356), .Z(n1396) );
  or2f U1160 ( .A1(n1400), .A2(n1401), .Z(n1352) );
  and2f U1176 ( .A1(n1414), .A2(n1415), .Z(c9) );
  and2f U1178 ( .A1(n1416), .A2(n1756), .Z(n1414) );
  or2f U1179 ( .A1(n1093), .A2(n1417), .Z(n1416) );
  or2f U1182 ( .A1(n1421), .A2(v3), .Z(n1420) );
  and2f U1185 ( .A1(n1423), .A2(n1424), .Z(n1422) );
  or2f U1195 ( .A1(b), .A2(n1432), .Z(n1431) );
  and2f U1196 ( .A1(n1433), .A2(n1193), .Z(n1432) );
  or2f U1197 ( .A1(n1434), .A2(n1435), .Z(n1433) );
  or2f U1202 ( .A1(n1438), .A2(n1401), .Z(n1437) );
  or2f U1203 ( .A1(n1439), .A2(n285), .Z(n1401) );
  inv1f U1252 ( .I(n1473), .ZN(n1167) );
  or2f U1254 ( .A1(n1474), .A2(f0), .Z(n1473) );
  and2f U1255 ( .A1(n1475), .A2(n1476), .Z(n1474) );
  and2f U1258 ( .A1(n1481), .A2(s4), .Z(n1475) );
  or2f U1263 ( .A1(n1486), .A2(q5), .Z(n1484) );
  inv1f U1264 ( .I(n1487), .ZN(n1486) );
  or2f U1265 ( .A1(n1488), .A2(n1489), .Z(n1487) );
  or2f U1266 ( .A1(x4), .A2(y4), .Z(n1489) );
  or2f U1267 ( .A1(n1955), .A2(w4), .Z(n1488) );
  or2f U1283 ( .A1(n1502), .A2(u1), .Z(n1501) );
  or2f U1285 ( .A1(n1503), .A2(n1504), .Z(n1502) );
  or2f U1304 ( .A1(n1520), .A2(n1521), .Z(n1519) );
  or2f U1305 ( .A1(n1522), .A2(n1523), .Z(n1521) );
  and2f U1325 ( .A1(n827), .A2(p4), .Z(n960) );
  and2f U1326 ( .A1(n959), .A2(g4), .Z(n827) );
  and2f U1331 ( .A1(d4), .A2(n1539), .Z(n986) );
  and2f U1332 ( .A1(e4), .A2(f4), .Z(n1539) );
  and2f U1333 ( .A1(q5), .A2(n1540), .Z(n1538) );
  and2f U1348 ( .A1(t3), .A2(n1551), .Z(n1548) );
  and2f U1351 ( .A1(n2038), .A2(n1534), .Z(n1554) );
  or2f U1355 ( .A1(n1751), .A2(n325), .Z(n260) );
  or2f U1359 ( .A1(n1556), .A2(h0), .Z(n410) );
  and2f U1360 ( .A1(n1557), .A2(p3), .Z(n1556) );
  or2f U1362 ( .A1(n1558), .A2(h0), .Z(n777) );
  and2f U1363 ( .A1(i3), .A2(n900), .Z(n1558) );
  and2f U1365 ( .A1(h3), .A2(n1561), .Z(n1560) );
  or2f U1366 ( .A1(n1562), .A2(n935), .Z(n1561) );
  or2f U1369 ( .A1(n1563), .A2(n402), .Z(n254) );
  or2f U1372 ( .A1(d0), .A2(n1566), .Z(n1565) );
  and2f U1389 ( .A1(n2038), .A2(n319), .Z(n1563) );
  or2f U1394 ( .A1(n562), .A2(p3), .Z(n1581) );
  and2f U1399 ( .A1(p5), .A2(n1585), .Z(n1559) );
  or2f U1416 ( .A1(n1591), .A2(n1018), .Z(a8) );
  and2f U1418 ( .A1(n261), .A2(n1592), .Z(n1591) );
  or2f U1419 ( .A1(n1593), .A2(n1594), .Z(n1592) );
  or2f U1421 ( .A1(n1596), .A2(t2), .Z(n1595) );
  and2f U1422 ( .A1(t2), .A2(n1596), .Z(n1593) );
  or2f U1423 ( .A1(n1597), .A2(n269), .Z(n1596) );
  inv1f U1424 ( .I(n333), .ZN(n269) );
  or2f U1426 ( .A1(f), .A2(n1600), .Z(n1599) );
  and2f U1436 ( .A1(n1609), .A2(n1610), .Z(n1597) );
  or2f U1437 ( .A1(n1611), .A2(n2023), .Z(n1610) );
  or2f U1440 ( .A1(n1612), .A2(n1613), .Z(n1387) );
  and2f U1441 ( .A1(s2), .A2(n1614), .Z(n1613) );
  or2f U1442 ( .A1(n1615), .A2(n273), .Z(n1614) );
  and2f U1447 ( .A1(n1617), .A2(n1618), .Z(n1390) );
  or2f U1450 ( .A1(n276), .A2(s2), .Z(n1617) );
  and2f U1451 ( .A1(n274), .A2(n1620), .Z(n276) );
  and2f U1454 ( .A1(n2065), .A2(n2041), .Z(n1615) );
  and2f U1455 ( .A1(n695), .A2(n2065), .Z(n1619) );
  and2f U1457 ( .A1(n699), .A2(m1), .Z(n1621) );
  and2f U1468 ( .A1(n1627), .A2(n1754), .Z(n1625) );
  or2f U1469 ( .A1(n1207), .A2(n1628), .Z(n1627) );
  or2f U1470 ( .A1(n1629), .A2(n1630), .Z(n1628) );
  or2f U1472 ( .A1(n1632), .A2(t1), .Z(n1631) );
  and2f U1475 ( .A1(n1634), .A2(n1635), .Z(n1633) );
  inv1f U1496 ( .I(n287), .ZN(n285) );
  or2f U1497 ( .A1(n1643), .A2(h), .Z(n287) );
  and2f U1498 ( .A1(n1644), .A2(n1645), .Z(n1643) );
  and2f U1504 ( .A1(n1647), .A2(w0), .Z(n1644) );
  inv1f U1526 ( .I(n1), .ZN(n699) );
  or2f U1604 ( .A1(n1957), .A2(n2050), .Z(n1715) );
  or2f U1610 ( .A1(n1993), .A2(n1718), .Z(n1717) );
  inv1f U1611 ( .I(o1), .ZN(n1718) );
  or2f U1614 ( .A1(n1722), .A2(n1723), .Z(n1721) );
  inv1f U1616 ( .I(o5), .ZN(n1723) );
  or2 U1618 ( .A1(n1925), .A2(n1815), .Z(n1725) );
  buf0 U1625 ( .I(a), .Z(l6) );
  buf0 U1626 ( .I(e1), .Z(m6) );
  buf0 U1627 ( .I(n1970), .Z(n6) );
  buf0 U1628 ( .I(j1), .Z(r6) );
  buf0 U1629 ( .I(n1969), .Z(v6) );
  buf0 U1630 ( .I(y), .Z(h10) );
  buf0 U1631 ( .I(a5), .Z(i10) );
  buf0 U1632 ( .I(n1968), .Z(j10) );
  buf0 U1633 ( .I(n1967), .Z(o10) );
  buf0 U1634 ( .I(g5), .Z(p10) );
  buf0 U1635 ( .I(n1966), .Z(v10) );
  or2f U1636 ( .A1(n1549), .A2(n1744), .Z(n1742) );
  and2f U1637 ( .A1(n1742), .A2(n1743), .Z(a9) );
  or2 U1638 ( .A1(n246), .A2(n247), .Z(n1743) );
  or2f U1639 ( .A1(n1548), .A2(n246), .Z(n1744) );
  or2f U1640 ( .A1(n260), .A2(n1747), .Z(n1745) );
  and2f U1641 ( .A1(n1745), .A2(n1746), .Z(n1552) );
  or2f U1643 ( .A1(n1554), .A2(n252), .Z(n1747) );
  inv1 U1646 ( .I(n1749), .ZN(n845) );
  and2 U1648 ( .A1(n259), .A2(n1751), .Z(n324) );
  and2 U1649 ( .A1(j5), .A2(n1749), .Z(n844) );
  and2 U1650 ( .A1(n751), .A2(n1749), .Z(n1846) );
  and2 U1651 ( .A1(r4), .A2(n1749), .Z(n1698) );
  and2 U1653 ( .A1(n321), .A2(n1730), .Z(n314) );
  or2 U1656 ( .A1(z), .A2(n1012), .Z(l9) );
  or2 U1657 ( .A1(z), .A2(n1016), .Z(k9) );
  or2 U1658 ( .A1(z), .A2(n1265), .Z(n1264) );
  or2 U1659 ( .A1(z), .A2(n1317), .Z(n1316) );
  or2 U1660 ( .A1(z), .A2(n1077), .Z(n1076) );
  or2 U1661 ( .A1(z), .A2(n1119), .Z(n1118) );
  or2 U1662 ( .A1(z), .A2(n1214), .Z(n1213) );
  or2 U1663 ( .A1(n845), .A2(n846), .Z(n842) );
  and2 U1664 ( .A1(j5), .A2(n845), .Z(n881) );
  or2 U1665 ( .A1(n845), .A2(n1936), .Z(n1937) );
  or2 U1666 ( .A1(n845), .A2(n1843), .Z(n1844) );
  or2 U1667 ( .A1(z), .A2(n961), .Z(n1690) );
  or2 U1668 ( .A1(n845), .A2(n1955), .Z(n1762) );
  or2f U1678 ( .A1(b5), .A2(n1757), .Z(n1931) );
  or2f U1680 ( .A1(n1721), .A2(i5), .Z(n1833) );
  inv1f U1681 ( .I(n1833), .ZN(n1823) );
  and2f U1682 ( .A1(n1931), .A2(n1823), .Z(n1759) );
  and2f U1683 ( .A1(n1936), .A2(n1833), .Z(n1758) );
  or2f U1684 ( .A1(n1759), .A2(n1758), .Z(n1763) );
  and2f U1685 ( .A1(n1936), .A2(n1763), .Z(n1760) );
  and2f U1686 ( .A1(n1835), .A2(n1760), .Z(n1761) );
  or2f U1687 ( .A1(n1761), .A2(e5), .Z(n1968) );
  inv1f U1694 ( .I(n1906), .ZN(n1901) );
  or2f U1698 ( .A1(n1901), .A2(n1767), .Z(n1905) );
  or2f U1723 ( .A1(n1717), .A2(k1), .Z(n1840) );
  inv1f U1724 ( .I(n1840), .ZN(n1837) );
  and2f U1725 ( .A1(n1886), .A2(n1837), .Z(n1779) );
  and2f U1726 ( .A1(n1879), .A2(n2028), .Z(n1778) );
  or2f U1727 ( .A1(n1779), .A2(n1778), .Z(n1785) );
  and2f U1728 ( .A1(n1879), .A2(n1785), .Z(n1780) );
  and2f U1729 ( .A1(n1842), .A2(n1780), .Z(n1781) );
  or2f U1730 ( .A1(n1781), .A2(i1), .Z(n1970) );
  or2f U1731 ( .A1(n1970), .A2(g1), .Z(n1786) );
  or2f U1735 ( .A1(n1986), .A2(n286), .Z(n1635) );
  or2f U1743 ( .A1(n1970), .A2(n2029), .Z(n1787) );
  or2f U1744 ( .A1(n1787), .A2(h1), .Z(n1804) );
  and2f U1745 ( .A1(n1969), .A2(n1804), .Z(n1788) );
  and2f U1746 ( .A1(n1789), .A2(n1788), .Z(n1600) );
  and2f U1754 ( .A1(n1793), .A2(n1966), .Z(n1794) );
  and2f U1760 ( .A1(n1300), .A2(n1819), .Z(n1439) );
  or2f U1762 ( .A1(n1797), .A2(g0), .Z(n1820) );
  inv1f U1764 ( .I(n1820), .ZN(n1821) );
  or2f U1772 ( .A1(n1799), .A2(n2036), .Z(n1854) );
  or2f U1776 ( .A1(n1849), .A2(n1801), .Z(n1853) );
  and2f U1790 ( .A1(n1173), .A2(n1821), .Z(n1324) );
  and2f U1792 ( .A1(n1295), .A2(n1819), .Z(n1294) );
  and2f U1805 ( .A1(z4), .A2(n1725), .Z(n1817) );
  or2f U1807 ( .A1(n1817), .A2(n1816), .Z(n1258) );
  and2f U1814 ( .A1(n1168), .A2(n1821), .Z(n1166) );
  and2f U1833 ( .A1(d1), .A2(n1720), .Z(n1831) );
  inv1f U1896 ( .I(n1889), .ZN(n1890) );
  or2f U1897 ( .A1(n1890), .A2(n1961), .Z(n1891) );
  and2f U1898 ( .A1(n1891), .A2(d1), .Z(n1892) );
  inv1f U1944 ( .I(n1940), .ZN(n1941) );
  or2f U1945 ( .A1(n1941), .A2(n1955), .Z(n1942) );
  and2f U1946 ( .A1(n1942), .A2(z4), .Z(n1943) );
  or2 U1609 ( .A1(n1302), .A2(n1303), .Z(n1301) );
  or2f U1612 ( .A1(n1205), .A2(n1206), .Z(n1203) );
  and2 U1613 ( .A1(n1203), .A2(n1818), .Z(n1200) );
  and2f U1615 ( .A1(n1506), .A2(n1986), .Z(n1505) );
  inv1f U1617 ( .I(n1981), .ZN(n695) );
  inv1f U1619 ( .I(n777), .ZN(n473) );
  inv1f U1620 ( .I(n960), .ZN(n1009) );
  inv1f U1621 ( .I(n982), .ZN(n981) );
  or2f U1622 ( .A1(n1853), .A2(n1719), .Z(n1866) );
  or2f U1623 ( .A1(n1293), .A2(n1250), .Z(n1292) );
  inv1f U1624 ( .I(n1931), .ZN(n1936) );
  or2f U1642 ( .A1(n1564), .A2(n1565), .Z(n2049) );
  or2f U1644 ( .A1(f1), .A2(n1777), .Z(n1886) );
  inv1f U1645 ( .I(n1886), .ZN(n1879) );
  and2 U1647 ( .A1(g3), .A2(n965), .Z(n966) );
  inv1 U1652 ( .I(n2060), .ZN(n2062) );
  or2 U1654 ( .A1(n1728), .A2(c5), .Z(n2005) );
  and2 U1655 ( .A1(n897), .A2(n898), .Z(n896) );
  inv1 U1669 ( .I(n1501), .ZN(n1500) );
  and2 U1670 ( .A1(u1), .A2(n1502), .Z(n1499) );
  and2 U1671 ( .A1(n1436), .A2(n1403), .Z(n1435) );
  inv1 U1672 ( .I(n1398), .ZN(n1397) );
  and2 U1673 ( .A1(n1291), .A2(n1252), .Z(n1290) );
  inv1 U1674 ( .I(n1292), .ZN(n1291) );
  and2 U1675 ( .A1(y1), .A2(n1292), .Z(n1289) );
  or2 U1676 ( .A1(n1284), .A2(n1183), .Z(n1341) );
  inv1 U1677 ( .I(n1280), .ZN(n1279) );
  or2 U1679 ( .A1(n1142), .A2(n1101), .Z(n1141) );
  inv1 U1688 ( .I(n1054), .ZN(n1053) );
  and2 U1689 ( .A1(n321), .A2(n777), .Z(n774) );
  or2 U1690 ( .A1(n609), .A2(n610), .Z(n608) );
  or2 U1691 ( .A1(n552), .A2(o3), .Z(n551) );
  or2 U1692 ( .A1(n468), .A2(n469), .Z(n467) );
  or2 U1693 ( .A1(n1925), .A2(n1924), .Z(n1927) );
  or2 U1695 ( .A1(n1831), .A2(n1830), .Z(n1065) );
  and2 U1696 ( .A1(n782), .A2(n783), .Z(n781) );
  or2 U1697 ( .A1(n574), .A2(y1), .Z(n782) );
  inv1 U1699 ( .I(n1022), .ZN(n1021) );
  or2 U1700 ( .A1(n965), .A2(g3), .Z(n964) );
  and2 U1701 ( .A1(h3), .A2(n929), .Z(n926) );
  and2 U1702 ( .A1(n665), .A2(n247), .Z(t8) );
  and2 U1703 ( .A1(n406), .A2(n407), .Z(n397) );
  and2 U1704 ( .A1(n311), .A2(n247), .Z(y8) );
  or2f U1705 ( .A1(n1991), .A2(n1992), .Z(n333) );
  inv1f U1706 ( .I(n1854), .ZN(n1849) );
  inv1f U1707 ( .I(n1818), .ZN(n1986) );
  and2 U1708 ( .A1(n274), .A2(n275), .Z(n271) );
  inv1 U1709 ( .I(n275), .ZN(n2023) );
  inv1 U1710 ( .I(n275), .ZN(n2022) );
  or2f U1711 ( .A1(n1784), .A2(g), .Z(n275) );
  or2f U1712 ( .A1(n1866), .A2(n1827), .Z(n1873) );
  or2f U1713 ( .A1(n1764), .A2(d5), .Z(n2012) );
  or2f U1714 ( .A1(y2), .A2(n1147), .Z(n1239) );
  and2f U1715 ( .A1(v1), .A2(n1819), .Z(n1400) );
  or2f U1716 ( .A1(n1973), .A2(n473), .Z(n558) );
  and2f U1717 ( .A1(n2063), .A2(n1586), .Z(n937) );
  and2 U1718 ( .A1(n2002), .A2(n2003), .Z(n1971) );
  inv1 U1719 ( .I(n259), .ZN(n2038) );
  or2f U1720 ( .A1(n1323), .A2(n1273), .Z(n1322) );
  and2f U1721 ( .A1(n410), .A2(q3), .Z(n1730) );
  inv1f U1722 ( .I(n1818), .ZN(n1819) );
  and2f U1732 ( .A1(n2009), .A2(n2010), .Z(n319) );
  and2 U1733 ( .A1(n2021), .A2(n2037), .Z(n780) );
  or2 U1734 ( .A1(n1165), .A2(n1127), .Z(n1164) );
  and2 U1736 ( .A1(n2038), .A2(n470), .Z(n469) );
  inv1 U1737 ( .I(j), .ZN(n1144) );
  inv1 U1738 ( .I(n1106), .ZN(n2046) );
  inv1 U1739 ( .I(n1108), .ZN(n1101) );
  or2 U1740 ( .A1(n2046), .A2(n2047), .Z(n2045) );
  or2 U1741 ( .A1(n560), .A2(n561), .Z(n559) );
  inv1 U1742 ( .I(n1730), .ZN(n1751) );
  or2 U1747 ( .A1(n1222), .A2(n1223), .Z(n1221) );
  or2 U1748 ( .A1(n1809), .A2(n1447), .Z(n1810) );
  or2 U1749 ( .A1(n1808), .A2(n1807), .Z(n1809) );
  or2 U1750 ( .A1(c), .A2(n1896), .Z(n2059) );
  and2 U1751 ( .A1(n835), .A2(n788), .Z(n834) );
  and2 U1752 ( .A1(m2), .A2(n572), .Z(n683) );
  or2 U1753 ( .A1(n521), .A2(n876), .Z(n566) );
  and2 U1755 ( .A1(n2037), .A2(n970), .Z(n969) );
  inv1 U1756 ( .I(n894), .ZN(n893) );
  or2 U1757 ( .A1(n779), .A2(n466), .Z(n778) );
  and2 U1758 ( .A1(n1974), .A2(n321), .Z(n668) );
  or2 U1759 ( .A1(n466), .A2(n612), .Z(n676) );
  and2 U1761 ( .A1(n2037), .A2(n560), .Z(n609) );
  inv1 U1763 ( .I(n464), .ZN(n463) );
  inv1 U1765 ( .I(n408), .ZN(n407) );
  and2 U1766 ( .A1(w3), .A2(n1371), .Z(n1368) );
  and2 U1767 ( .A1(n1163), .A2(n1129), .Z(n1162) );
  and2 U1768 ( .A1(n660), .A2(n602), .Z(n659) );
  and2 U1769 ( .A1(o4), .A2(n393), .Z(n543) );
  or2 U1770 ( .A1(n1905), .A2(n1959), .Z(n1912) );
  or2 U1771 ( .A1(n1912), .A2(n1958), .Z(n1914) );
  or2 U1773 ( .A1(n1773), .A2(n1690), .Z(n1774) );
  or2 U1774 ( .A1(n1772), .A2(n1692), .Z(n1773) );
  and2 U1775 ( .A1(g5), .A2(n981), .Z(n980) );
  and2 U1777 ( .A1(n1006), .A2(n1756), .Z(n1005) );
  or2 U1778 ( .A1(n2056), .A2(n1949), .Z(n2027) );
  or2 U1779 ( .A1(a0), .A2(n1946), .Z(n2056) );
  and2 U1780 ( .A1(n2006), .A2(n2007), .Z(n1582) );
  or2 U1781 ( .A1(h3), .A2(i3), .Z(n2008) );
  and2 U1782 ( .A1(n1301), .A2(n1297), .Z(n1251) );
  and2 U1783 ( .A1(q2), .A2(r2), .Z(n273) );
  inv1 U1784 ( .I(q5), .ZN(n2064) );
  inv1 U1785 ( .I(n1559), .ZN(n1584) );
  or2 U1786 ( .A1(n1559), .A2(n1560), .Z(n900) );
  inv1 U1787 ( .I(j1), .ZN(n1993) );
  inv1 U1788 ( .I(r1), .ZN(n1961) );
  or2 U1789 ( .A1(n1401), .A2(n1995), .Z(n1398) );
  and2 U1791 ( .A1(n1389), .A2(n1144), .Z(n1147) );
  inv1 U1793 ( .I(n1138), .ZN(n1137) );
  and2 U1794 ( .A1(n1143), .A2(n1144), .Z(n1139) );
  or2 U1795 ( .A1(n1145), .A2(n1146), .Z(n1143) );
  inv1 U1796 ( .I(n2014), .ZN(n1566) );
  inv1 U1797 ( .I(n2013), .ZN(n2015) );
  and2 U1798 ( .A1(n1583), .A2(n1584), .Z(n901) );
  or2 U1799 ( .A1(n937), .A2(h3), .Z(n1583) );
  or2 U1800 ( .A1(n2021), .A2(n1971), .Z(n472) );
  inv1 U1801 ( .I(n404), .ZN(n403) );
  or2 U1802 ( .A1(n1581), .A2(n470), .Z(n1579) );
  inv1 U1803 ( .I(n259), .ZN(n2037) );
  or2 U1804 ( .A1(n470), .A2(q3), .Z(n2011) );
  inv1 U1806 ( .I(j0), .ZN(n1540) );
  or2 U1808 ( .A1(z), .A2(n1957), .Z(n746) );
  inv1 U1809 ( .I(l5), .ZN(n1957) );
  and2 U1810 ( .A1(n1785), .A2(n1727), .Z(n1726) );
  or2 U1811 ( .A1(n1717), .A2(k1), .Z(n2028) );
  inv1 U1812 ( .I(e1), .ZN(n1777) );
  and2 U1813 ( .A1(t1), .A2(n1632), .Z(n1629) );
  inv1 U1815 ( .I(n1631), .ZN(n1630) );
  and2 U1816 ( .A1(v1), .A2(n1437), .Z(n1434) );
  inv1 U1817 ( .I(n1437), .ZN(n1436) );
  and2 U1818 ( .A1(x1), .A2(n1351), .Z(n1348) );
  and2 U1819 ( .A1(z1), .A2(n1247), .Z(n1244) );
  and2 U1820 ( .A1(a2), .A2(n1197), .Z(n1194) );
  inv1 U1821 ( .I(n1196), .ZN(n1195) );
  and2 U1822 ( .A1(q1), .A2(n1040), .Z(n1038) );
  inv1 U1823 ( .I(l), .ZN(n1040) );
  inv1 U1824 ( .I(n1595), .ZN(n1594) );
  inv1 U1825 ( .I(n1185), .ZN(n1184) );
  or2 U1826 ( .A1(n1105), .A2(n1058), .Z(n1104) );
  or2 U1827 ( .A1(n324), .A2(n325), .Z(n323) );
  and2 U1828 ( .A1(z3), .A2(n1219), .Z(n1216) );
  inv1 U1829 ( .I(n1219), .ZN(n1218) );
  inv1 U1830 ( .I(n1082), .ZN(n1081) );
  and2 U1831 ( .A1(n889), .A2(i4), .Z(n888) );
  or2 U1832 ( .A1(n1538), .A2(n986), .Z(n889) );
  inv1 U1834 ( .I(n390), .ZN(n389) );
  or2 U1835 ( .A1(n2019), .A2(n393), .Z(n390) );
  or2 U1836 ( .A1(n1765), .A2(n2012), .Z(n1906) );
  inv1 U1837 ( .I(n1762), .ZN(n1765) );
  and2 U1838 ( .A1(n1763), .A2(n1729), .Z(n1728) );
  inv1 U1839 ( .I(g5), .ZN(n1722) );
  or2 U1840 ( .A1(z), .A2(n1001), .Z(n1000) );
  inv1 U1841 ( .I(n1002), .ZN(n1001) );
  or2 U1842 ( .A1(n1003), .A2(n981), .Z(n1002) );
  inv1 U1843 ( .I(a5), .ZN(n1757) );
  or2 U1844 ( .A1(n498), .A2(n499), .Z(w5) );
  or2 U1845 ( .A1(n508), .A2(n509), .Z(n498) );
  or2 U1846 ( .A1(n1508), .A2(n1509), .Z(b6) );
  or2 U1847 ( .A1(n1518), .A2(n1519), .Z(n1508) );
  or2 U1848 ( .A1(n1858), .A2(y0), .Z(n1859) );
  and2 U1849 ( .A1(n1951), .A2(n1871), .Z(n1874) );
  and2 U1850 ( .A1(n1951), .A2(n1720), .Z(n1878) );
  inv1 U1851 ( .I(n1875), .ZN(n1876) );
  and2 U1852 ( .A1(n1951), .A2(n1065), .Z(k6) );
  and2 U1853 ( .A1(n1890), .A2(n1068), .Z(n1830) );
  and2 U1854 ( .A1(n1900), .A2(n1754), .Z(t6) );
  and2 U1855 ( .A1(n282), .A2(n1498), .Z(n1496) );
  or2 U1856 ( .A1(n1499), .A2(n1500), .Z(n1498) );
  or2 U1857 ( .A1(n1391), .A2(n1392), .Z(d7) );
  and2 U1858 ( .A1(n282), .A2(n1288), .Z(n1286) );
  or2 U1859 ( .A1(n1289), .A2(n1290), .Z(n1288) );
  and2 U1860 ( .A1(n834), .A2(n574), .Z(n833) );
  or2 U1861 ( .A1(n679), .A2(b), .Z(t7) );
  and2 U1862 ( .A1(n680), .A2(n681), .Z(n679) );
  and2 U1863 ( .A1(n327), .A2(n261), .Z(y7) );
  inv1 U1864 ( .I(n265), .ZN(n264) );
  or2 U1865 ( .A1(n1183), .A2(n1383), .Z(n1378) );
  or2 U1866 ( .A1(n1340), .A2(n1341), .Z(n1331) );
  and2 U1867 ( .A1(n261), .A2(n1276), .Z(f8) );
  or2 U1868 ( .A1(n1277), .A2(n1278), .Z(n1276) );
  and2 U1869 ( .A1(z2), .A2(n1231), .Z(n1228) );
  and2 U1870 ( .A1(n1140), .A2(n1141), .Z(n1132) );
  and2 U1871 ( .A1(e3), .A2(n1023), .Z(n1020) );
  and2 U1872 ( .A1(n963), .A2(n964), .Z(n962) );
  inv1 U1873 ( .I(n966), .ZN(n963) );
  and2 U1874 ( .A1(n247), .A2(n925), .Z(o8) );
  inv1 U1875 ( .I(n928), .ZN(n927) );
  or2 U1876 ( .A1(n890), .A2(n246), .Z(p8) );
  and2 U1877 ( .A1(i3), .A2(n895), .Z(n892) );
  and2 U1878 ( .A1(n771), .A2(n247), .Z(s8) );
  or2 U1879 ( .A1(n673), .A2(n778), .Z(n772) );
  or2 U1880 ( .A1(n675), .A2(n676), .Z(n666) );
  and2 U1881 ( .A1(n247), .A2(n603), .Z(u8) );
  or2 U1882 ( .A1(n604), .A2(n605), .Z(n603) );
  and2 U1883 ( .A1(n3), .A2(n607), .Z(n604) );
  inv1 U1884 ( .I(n551), .ZN(n550) );
  and2 U1885 ( .A1(p3), .A2(n465), .Z(n462) );
  or2 U1886 ( .A1(n395), .A2(n246), .Z(x8) );
  and2 U1887 ( .A1(s3), .A2(n253), .Z(n249) );
  inv1 U1888 ( .I(n1550), .ZN(n1549) );
  or2 U1889 ( .A1(n1079), .A2(m3), .Z(n1415) );
  and2 U1890 ( .A1(n1159), .A2(n1367), .Z(n1365) );
  or2 U1891 ( .A1(n1315), .A2(n1316), .Z(e9) );
  and2 U1892 ( .A1(n1318), .A2(n1079), .Z(n1317) );
  and2 U1893 ( .A1(n1159), .A2(n1160), .Z(n1156) );
  or2 U1894 ( .A1(n1161), .A2(n1162), .Z(n1160) );
  and2 U1895 ( .A1(n659), .A2(n394), .Z(n658) );
  or2 U1899 ( .A1(n539), .A2(z), .Z(v9) );
  and2 U1900 ( .A1(n540), .A2(n541), .Z(n539) );
  or2 U1901 ( .A1(n1910), .A2(u4), .Z(n1911) );
  and2 U1902 ( .A1(n1954), .A2(n1923), .Z(n1926) );
  and2 U1903 ( .A1(n1954), .A2(n1258), .Z(g10) );
  and2 U1904 ( .A1(n1941), .A2(n1261), .Z(n1816) );
  or2 U1905 ( .A1(n979), .A2(n980), .Z(n978) );
  and2 U1906 ( .A1(n1950), .A2(n1756), .Z(t10) );
  and2 U1907 ( .A1(n2025), .A2(n2026), .Z(n1950) );
  inv1f U1908 ( .I(h0), .ZN(n1580) );
  and2 U1909 ( .A1(n2063), .A2(n1971), .Z(n933) );
  inv1 U1910 ( .I(n320), .ZN(n1972) );
  inv1 U1911 ( .I(n320), .ZN(n402) );
  or2 U1912 ( .A1(n896), .A2(n1972), .Z(n895) );
  and2 U1913 ( .A1(n1972), .A2(s0), .Z(n1522) );
  inv1 U1914 ( .I(n2063), .ZN(n1562) );
  and2 U1915 ( .A1(n1750), .A2(m5), .Z(n1749) );
  or2 U1916 ( .A1(n612), .A2(n673), .Z(n1973) );
  and2 U1917 ( .A1(n777), .A2(l3), .Z(n1974) );
  inv1 U1918 ( .I(n1974), .ZN(n611) );
  or2f U1919 ( .A1(n550), .A2(n1977), .Z(n1975) );
  and2 U1920 ( .A1(n1975), .A2(n1976), .Z(v8) );
  or2 U1921 ( .A1(n246), .A2(n247), .Z(n1976) );
  or2f U1922 ( .A1(n549), .A2(n246), .Z(n1977) );
  and2 U1923 ( .A1(b4), .A2(n1821), .Z(n1087) );
  and2 U1924 ( .A1(y3), .A2(n1821), .Z(n1223) );
  and2 U1925 ( .A1(x3), .A2(n1821), .Z(n1272) );
  and2 U1926 ( .A1(a4), .A2(n1821), .Z(n1126) );
  or2 U1927 ( .A1(n1821), .A2(n1425), .Z(n1424) );
  and2 U1928 ( .A1(n2068), .A2(n1612), .Z(n1983) );
  inv1 U1929 ( .I(n1612), .ZN(n1618) );
  and2f U1930 ( .A1(p1), .A2(n1619), .Z(n1612) );
  and2 U1931 ( .A1(n1151), .A2(v2), .Z(n1188) );
  or2f U1932 ( .A1(n1402), .A2(n1403), .Z(n1357) );
  or2 U1933 ( .A1(n1784), .A2(g), .Z(n1978) );
  and2 U1934 ( .A1(n2022), .A2(n705), .Z(n1027) );
  inv1f U1935 ( .I(r5), .ZN(n1955) );
  or2 U1936 ( .A1(n1167), .A2(n1374), .Z(n1373) );
  or2 U1937 ( .A1(n1167), .A2(n1422), .Z(n1421) );
  and2 U1938 ( .A1(n2022), .A2(n1237), .Z(n1232) );
  and2 U1939 ( .A1(n2022), .A2(n1238), .Z(n1282) );
  and2 U1940 ( .A1(n1235), .A2(n275), .Z(n1234) );
  or2f U1941 ( .A1(n1598), .A2(n1599), .Z(n1979) );
  and2 U1942 ( .A1(q1), .A2(l1), .Z(n1980) );
  or2 U1943 ( .A1(b), .A2(n1775), .Z(n1981) );
  and2 U1947 ( .A1(n1614), .A2(n1984), .Z(n1982) );
  or2f U1948 ( .A1(n1982), .A2(n1983), .Z(n2066) );
  and2 U1949 ( .A1(s2), .A2(n2068), .Z(n1984) );
  or2f U1950 ( .A1(n1968), .A2(n2005), .Z(n1764) );
  and2 U1951 ( .A1(n1978), .A2(n1236), .Z(n1283) );
  or2f U1952 ( .A1(n1978), .A2(u2), .Z(n1187) );
  and2 U1953 ( .A1(n1621), .A2(n695), .Z(n1953) );
  inv1 U1954 ( .I(n1986), .ZN(n1985) );
  and2 U1955 ( .A1(z1), .A2(n1819), .Z(n1201) );
  and2 U1956 ( .A1(w1), .A2(n1819), .Z(n1355) );
  or2f U1957 ( .A1(n1274), .A2(n1275), .Z(n1225) );
  and2f U1958 ( .A1(n556), .A2(n1971), .Z(n555) );
  and2f U1959 ( .A1(n1650), .A2(n1825), .Z(n1649) );
  and2f U1960 ( .A1(n1102), .A2(n1151), .Z(n1380) );
  and2f U1961 ( .A1(n1102), .A2(n1103), .Z(n1097) );
  or2 U1962 ( .A1(n1853), .A2(n1987), .Z(n1889) );
  or2 U1963 ( .A1(n1719), .A2(n2057), .Z(n1987) );
  or2f U1964 ( .A1(n1892), .A2(n1990), .Z(n1988) );
  and2 U1965 ( .A1(n1988), .A2(n1989), .Z(n1900) );
  or2 U1966 ( .A1(n1899), .A2(n2058), .Z(n1989) );
  or2 U1967 ( .A1(n2059), .A2(n1899), .Z(n1990) );
  and2f U1968 ( .A1(n1788), .A2(n1789), .Z(n1991) );
  or2 U1969 ( .A1(n1598), .A2(f), .Z(n1992) );
  and2 U1970 ( .A1(d3), .A2(n1054), .Z(n1051) );
  and2f U1971 ( .A1(t2), .A2(n1387), .Z(n1386) );
  or2 U1972 ( .A1(n473), .A2(n474), .Z(n471) );
  inv1 U1973 ( .I(j1), .ZN(n479) );
  inv1 U1974 ( .I(n1996), .ZN(n1994) );
  or2f U1975 ( .A1(n1400), .A2(n1399), .Z(n1995) );
  and2 U1976 ( .A1(w1), .A2(n1398), .Z(n1395) );
  inv1 U1977 ( .I(n287), .ZN(n1996) );
  or2 U1978 ( .A1(n1996), .A2(n1505), .Z(n1504) );
  and2f U1979 ( .A1(n1561), .A2(n1999), .Z(n1997) );
  or2f U1980 ( .A1(n1997), .A2(n1998), .Z(n2051) );
  and2 U1981 ( .A1(n2053), .A2(n1559), .Z(n1998) );
  and2 U1982 ( .A1(h3), .A2(n2053), .Z(n1999) );
  and2f U1983 ( .A1(n1760), .A2(n1835), .Z(n2000) );
  or2f U1984 ( .A1(n2000), .A2(n2001), .Z(n1797) );
  or2 U1985 ( .A1(c5), .A2(e5), .Z(n2001) );
  or2 U1986 ( .A1(n2000), .A2(n2004), .Z(n2002) );
  and2f U1987 ( .A1(n2002), .A2(n2003), .Z(n259) );
  or2 U1988 ( .A1(e0), .A2(n1966), .Z(n2003) );
  or2 U1989 ( .A1(n2001), .A2(e0), .Z(n2004) );
  and2f U1990 ( .A1(n1969), .A2(n1786), .Z(n1784) );
  or2 U1991 ( .A1(n1551), .A2(t3), .Z(n1550) );
  and2 U1992 ( .A1(n1582), .A2(n1580), .Z(n562) );
  and2 U1993 ( .A1(n1579), .A2(n1580), .Z(n405) );
  and2 U1994 ( .A1(n259), .A2(n558), .Z(n610) );
  and2f U1995 ( .A1(n2043), .A2(n2023), .Z(n1100) );
  or2f U1996 ( .A1(n1905), .A2(n1724), .Z(n1918) );
  or2f U1997 ( .A1(n937), .A2(n2008), .Z(n2006) );
  or2 U1998 ( .A1(i3), .A2(n1584), .Z(n2007) );
  or2f U1999 ( .A1(n1581), .A2(n2011), .Z(n2009) );
  or2 U2000 ( .A1(q3), .A2(n1580), .Z(n2010) );
  and2 U2001 ( .A1(n1795), .A2(n1966), .Z(n2013) );
  or2f U2002 ( .A1(n1771), .A2(n2015), .Z(n2014) );
  or2f U2003 ( .A1(n1770), .A2(z), .Z(n1966) );
  or2 U2004 ( .A1(n1764), .A2(d5), .Z(n1793) );
  or2f U2005 ( .A1(n1918), .A2(n1813), .Z(n1925) );
  or2f U2006 ( .A1(n1786), .A2(i), .Z(n1818) );
  or2f U2007 ( .A1(n1961), .A2(a1), .Z(n1654) );
  or2f U2008 ( .A1(n986), .A2(n2018), .Z(n2016) );
  and2f U2009 ( .A1(n2016), .A2(n2017), .Z(n959) );
  or2 U2010 ( .A1(n1537), .A2(i4), .Z(n2017) );
  or2f U2011 ( .A1(n1538), .A2(n1537), .Z(n2018) );
  or2 U2012 ( .A1(n392), .A2(q4), .Z(n2019) );
  and2 U2013 ( .A1(n545), .A2(n392), .Z(n544) );
  and2 U2014 ( .A1(l2), .A2(k2), .Z(n2020) );
  and2 U2015 ( .A1(n685), .A2(n573), .Z(n684) );
  and2 U2016 ( .A1(n1582), .A2(n1580), .Z(n2021) );
  and2 U2017 ( .A1(n409), .A2(n319), .Z(n408) );
  inv1 U2018 ( .I(n319), .ZN(n318) );
  or2 U2019 ( .A1(n3), .A2(n2021), .Z(n561) );
  or2 U2020 ( .A1(n2022), .A2(b3), .Z(n1148) );
  or2 U2021 ( .A1(n2054), .A2(n1724), .Z(n2024) );
  or2f U2022 ( .A1(n1943), .A2(n2027), .Z(n2025) );
  or2 U2023 ( .A1(n1949), .A2(n2055), .Z(n2026) );
  and2f U2024 ( .A1(n259), .A2(n2049), .Z(n321) );
  or2 U2025 ( .A1(n1726), .A2(g1), .Z(n2029) );
  or2f U2026 ( .A1(n1390), .A2(n2032), .Z(n2030) );
  and2f U2027 ( .A1(n2030), .A2(n2031), .Z(n1145) );
  or2 U2028 ( .A1(a3), .A2(n1144), .Z(n2031) );
  or2 U2029 ( .A1(t2), .A2(a3), .Z(n2032) );
  or2f U2030 ( .A1(n1145), .A2(n2035), .Z(n2033) );
  and2f U2031 ( .A1(n2033), .A2(n2034), .Z(n1108) );
  or2 U2032 ( .A1(b3), .A2(n1144), .Z(n2034) );
  or2 U2033 ( .A1(n1146), .A2(b3), .Z(n2035) );
  or2f U2034 ( .A1(n1787), .A2(h1), .Z(n2036) );
  and2 U2035 ( .A1(n405), .A2(n2037), .Z(n400) );
  and2 U2036 ( .A1(n2038), .A2(n559), .Z(n553) );
  or2 U2037 ( .A1(n1554), .A2(n259), .Z(n1746) );
  and2f U2038 ( .A1(n2049), .A2(n2038), .Z(n317) );
  and2 U2039 ( .A1(r3), .A2(n2037), .Z(n257) );
  or2 U2040 ( .A1(n2038), .A2(n410), .Z(n404) );
  and2f U2041 ( .A1(n1794), .A2(n1795), .Z(n2039) );
  or2f U2042 ( .A1(n2039), .A2(n2040), .Z(n320) );
  or2 U2043 ( .A1(n1564), .A2(d0), .Z(n2040) );
  and2f U2044 ( .A1(n1980), .A2(n1754), .Z(n2041) );
  or2 U2045 ( .A1(n1058), .A2(n2047), .Z(n2042) );
  inv1 U2046 ( .I(b3), .ZN(n2047) );
  and2 U2047 ( .A1(q1), .A2(n1619), .Z(n2044) );
  and2 U2048 ( .A1(n1978), .A2(n2045), .Z(n1105) );
  or2f U2049 ( .A1(n1598), .A2(n1599), .Z(n2043) );
  inv1 U2050 ( .I(n2045), .ZN(n1103) );
  and2 U2051 ( .A1(n1978), .A2(n1979), .Z(n1102) );
  and2 U2052 ( .A1(n1138), .A2(n1979), .Z(n1140) );
  and2 U2053 ( .A1(n332), .A2(n1979), .Z(n330) );
  inv1 U2054 ( .I(n2044), .ZN(n274) );
  or2f U2055 ( .A1(n1564), .A2(n1565), .Z(n2048) );
  and2f U2056 ( .A1(n1329), .A2(w3), .Z(n1328) );
  and2f U2057 ( .A1(u3), .A2(v3), .Z(n1329) );
  or2f U2058 ( .A1(n1128), .A2(n1129), .Z(n1092) );
  and2f U2059 ( .A1(n1174), .A2(n1170), .Z(n1128) );
  and2 U2060 ( .A1(n967), .A2(n2048), .Z(n965) );
  and2 U2061 ( .A1(n404), .A2(n2048), .Z(n406) );
  and2 U2062 ( .A1(n672), .A2(n2048), .Z(n776) );
  and2f U2063 ( .A1(n1444), .A2(u1), .Z(n1443) );
  and2f U2064 ( .A1(s1), .A2(t1), .Z(n1444) );
  or2f U2065 ( .A1(n1251), .A2(n1252), .Z(n1206) );
  or2 U2066 ( .A1(n1024), .A2(n1104), .Z(n1095) );
  or2 U2067 ( .A1(n269), .A2(n336), .Z(n413) );
  and2 U2068 ( .A1(u), .A2(n269), .Z(n512) );
  or2 U2069 ( .A1(n269), .A2(n270), .Z(n268) );
  or2 U2070 ( .A1(n269), .A2(n1137), .Z(n1136) );
  or2f U2071 ( .A1(z), .A2(n5), .Z(n2050) );
  or2f U2072 ( .A1(n2051), .A2(n2052), .Z(n1557) );
  and2 U2073 ( .A1(k3), .A2(h0), .Z(n2052) );
  and2 U2074 ( .A1(i3), .A2(k3), .Z(n2053) );
  or2f U2075 ( .A1(n1552), .A2(n254), .Z(n1551) );
  or2 U2076 ( .A1(n254), .A2(n323), .Z(n312) );
  or2 U2077 ( .A1(n1972), .A2(n970), .Z(n990) );
  or2 U2078 ( .A1(n1972), .A2(n932), .Z(n931) );
  or2 U2079 ( .A1(n402), .A2(n403), .Z(n401) );
  or2f U2080 ( .A1(n2024), .A2(n1905), .Z(n1940) );
  or2 U2081 ( .A1(n1813), .A2(n1815), .Z(n2054) );
  or2 U2082 ( .A1(n1946), .A2(n1966), .Z(n2055) );
  or2 U2083 ( .A1(n1827), .A2(n1829), .Z(n2057) );
  or2 U2084 ( .A1(n1896), .A2(n1969), .Z(n2058) );
  or2 U2085 ( .A1(n1873), .A2(n1829), .Z(n1720) );
  inv1 U2086 ( .I(n1873), .ZN(n1870) );
  or2 U2087 ( .A1(n1873), .A2(n1872), .Z(n1875) );
  and2f U2088 ( .A1(n1580), .A2(m5), .Z(n2060) );
  or2f U2089 ( .A1(n1715), .A2(n2062), .Z(n2061) );
  inv1 U2090 ( .I(n2061), .ZN(n1585) );
  or2f U2091 ( .A1(n2064), .A2(n2061), .Z(n2063) );
  inv1 U2092 ( .I(n1715), .ZN(n1750) );
  and2f U2093 ( .A1(n1621), .A2(n1144), .Z(n2065) );
  or2f U2094 ( .A1(n2066), .A2(n2067), .Z(n1150) );
  and2 U2095 ( .A1(a3), .A2(j), .Z(n2067) );
  and2 U2096 ( .A1(t2), .A2(a3), .Z(n2068) );
  and2 U2097 ( .A1(n1169), .A2(n1170), .Z(n1168) );
  or2 U2098 ( .A1(n1171), .A2(n1172), .Z(n1169) );
  inv1 U2099 ( .I(y0), .ZN(n1963) );
  inv1 U2100 ( .I(x0), .ZN(n1964) );
  or2 U2101 ( .A1(n1965), .A2(n1800), .Z(n1801) );
  inv1 U2102 ( .I(w0), .ZN(n1800) );
  or2 U2103 ( .A1(n1960), .A2(n1766), .Z(n1767) );
  inv1 U2104 ( .I(s4), .ZN(n1766) );
  and2 U2105 ( .A1(n1296), .A2(n1297), .Z(n1295) );
  or2 U2106 ( .A1(n1298), .A2(n1299), .Z(n1296) );
  inv1 U2107 ( .I(n1894), .ZN(n1895) );
  and2 U2108 ( .A1(n1477), .A2(n1960), .Z(n1476) );
  inv1 U2109 ( .I(x3), .ZN(n1275) );
  inv1 U2110 ( .I(a4), .ZN(n1129) );
  inv1 U2111 ( .I(n1011), .ZN(n961) );
  inv1 U2112 ( .I(n748), .ZN(n538) );
  or2 U2113 ( .A1(n749), .A2(n750), .Z(n748) );
  or2 U2114 ( .A1(z), .A2(m5), .Z(n749) );
  or2 U2115 ( .A1(l5), .A2(n747), .Z(n750) );
  or2 U2116 ( .A1(n1826), .A2(n1964), .Z(n1719) );
  or2 U2117 ( .A1(n1963), .A2(n1825), .Z(n1826) );
  inv1 U2118 ( .I(q2), .ZN(n336) );
  and2 U2119 ( .A1(n1953), .A2(n1608), .Z(n1598) );
  or2 U2120 ( .A1(v0), .A2(n1961), .Z(n1608) );
  inv1 U2121 ( .I(f3), .ZN(n970) );
  and2 U2122 ( .A1(n1577), .A2(k5), .Z(n1564) );
  and2 U2123 ( .A1(n1578), .A2(n883), .Z(n1577) );
  or2 U2124 ( .A1(n1812), .A2(n1959), .Z(n1724) );
  or2 U2125 ( .A1(n1958), .A2(n1811), .Z(n1812) );
  or2 U2126 ( .A1(n648), .A2(n1952), .Z(n1946) );
  inv1 U2127 ( .I(k), .ZN(n1297) );
  inv1 U2128 ( .I(i0), .ZN(n1170) );
  or2 U2129 ( .A1(s1), .A2(t1), .Z(n1506) );
  and2 U2130 ( .A1(n1442), .A2(n1297), .Z(n1402) );
  inv1 U2131 ( .I(n1443), .ZN(n1442) );
  or2 U2132 ( .A1(n1356), .A2(n1357), .Z(n1302) );
  and2 U2133 ( .A1(y1), .A2(n1986), .Z(n1249) );
  and2 U2134 ( .A1(f3), .A2(g3), .Z(n935) );
  and2 U2135 ( .A1(n1375), .A2(n1821), .Z(n1374) );
  or2 U2136 ( .A1(u3), .A2(v3), .Z(n1375) );
  and2 U2137 ( .A1(n1327), .A2(n1170), .Z(n1274) );
  inv1 U2138 ( .I(n1328), .ZN(n1327) );
  or2 U2139 ( .A1(n1224), .A2(n1225), .Z(n1175) );
  or2 U2140 ( .A1(n1175), .A2(n1176), .Z(n1174) );
  or2 U2141 ( .A1(n1091), .A2(n1092), .Z(n1089) );
  inv1 U2142 ( .I(h5), .ZN(n1004) );
  inv1 U2143 ( .I(b1), .ZN(n1872) );
  or2 U2144 ( .A1(n1872), .A2(n1828), .Z(n1829) );
  inv1 U2145 ( .I(c1), .ZN(n1828) );
  inv1 U2146 ( .I(i1), .ZN(n1727) );
  or2 U2147 ( .A1(n1783), .A2(n1782), .Z(n1894) );
  or2 U2148 ( .A1(l1), .A2(n1), .Z(n1783) );
  or2 U2149 ( .A1(n1962), .A2(b), .Z(n1782) );
  and2 U2150 ( .A1(e3), .A2(n794), .Z(n520) );
  and2 U2151 ( .A1(c3), .A2(d3), .Z(n794) );
  and2 U2152 ( .A1(n699), .A2(n1962), .Z(n1657) );
  inv1 U2153 ( .I(n696), .ZN(n497) );
  or2 U2154 ( .A1(n697), .A2(n698), .Z(n696) );
  or2 U2155 ( .A1(m1), .A2(l1), .Z(n697) );
  or2 U2156 ( .A1(b), .A2(n699), .Z(n698) );
  inv1 U2157 ( .I(s1), .ZN(n286) );
  and2 U2158 ( .A1(n1646), .A2(n1965), .Z(n1645) );
  inv1 U2159 ( .I(v1), .ZN(n1403) );
  inv1 U2160 ( .I(w1), .ZN(n1356) );
  inv1 U2161 ( .I(y1), .ZN(n1252) );
  inv1 U2162 ( .I(z1), .ZN(n1205) );
  inv1 U2163 ( .I(n1661), .ZN(n1603) );
  or2 U2164 ( .A1(n1662), .A2(n1663), .Z(n1661) );
  or2 U2165 ( .A1(n1666), .A2(n1667), .Z(n1662) );
  or2 U2166 ( .A1(n1664), .A2(n1665), .Z(n1663) );
  and2 U2167 ( .A1(n909), .A2(n2), .Z(n521) );
  inv1 U2168 ( .I(n521), .ZN(n480) );
  or2 U2169 ( .A1(r2), .A2(q2), .Z(n1620) );
  inv1 U2170 ( .I(n273), .ZN(n272) );
  inv1 U2171 ( .I(n1387), .ZN(n1611) );
  inv1 U2172 ( .I(w2), .ZN(n1338) );
  inv1 U2173 ( .I(n1147), .ZN(n1337) );
  or2 U2174 ( .A1(w2), .A2(x2), .Z(n1238) );
  inv1 U2175 ( .I(u2), .ZN(n1146) );
  or2 U2176 ( .A1(g3), .A2(f3), .Z(n1586) );
  inv1 U2177 ( .I(n935), .ZN(n934) );
  inv1 U2178 ( .I(n900), .ZN(n899) );
  or2 U2179 ( .A1(n1820), .A2(u3), .Z(n1423) );
  inv1 U2180 ( .I(y3), .ZN(n1224) );
  inv1 U2181 ( .I(b4), .ZN(n1091) );
  inv1 U2182 ( .I(r4), .ZN(n1960) );
  inv1 U2183 ( .I(u4), .ZN(n1958) );
  inv1 U2184 ( .I(t4), .ZN(n1959) );
  inv1 U2185 ( .I(x4), .ZN(n1924) );
  inv1 U2186 ( .I(e5), .ZN(n1729) );
  and2 U2187 ( .A1(n1011), .A2(n1756), .Z(n1047) );
  inv1 U2188 ( .I(n5), .ZN(n747) );
  or2 U2189 ( .A1(n801), .A2(n802), .Z(n797) );
  and2 U2190 ( .A1(x1), .A2(q), .Z(n801) );
  or2 U2191 ( .A1(n803), .A2(n804), .Z(n802) );
  and2 U2192 ( .A1(t2), .A2(o), .Z(n803) );
  or2 U2193 ( .A1(n799), .A2(n800), .Z(n798) );
  and2 U2194 ( .A1(u1), .A2(r), .Z(n799) );
  and2 U2195 ( .A1(y0), .A2(w), .Z(n800) );
  or2 U2196 ( .A1(n807), .A2(n808), .Z(n806) );
  and2 U2197 ( .A1(j2), .A2(t), .Z(n807) );
  or2 U2198 ( .A1(n809), .A2(n810), .Z(n808) );
  and2 U2199 ( .A1(m), .A2(e3), .Z(n809) );
  or2 U2200 ( .A1(n811), .A2(n812), .Z(n805) );
  and2 U2201 ( .A1(d1), .A2(v), .Z(n811) );
  or2 U2202 ( .A1(n813), .A2(n814), .Z(n812) );
  and2 U2203 ( .A1(a2), .A2(p), .Z(n813) );
  or2 U2204 ( .A1(n722), .A2(n723), .Z(n718) );
  and2 U2205 ( .A1(w1), .A2(q), .Z(n722) );
  or2 U2206 ( .A1(n724), .A2(n725), .Z(n723) );
  and2 U2207 ( .A1(o), .A2(s2), .Z(n724) );
  or2 U2208 ( .A1(n720), .A2(n721), .Z(n719) );
  and2 U2209 ( .A1(t1), .A2(r), .Z(n720) );
  and2 U2210 ( .A1(x0), .A2(w), .Z(n721) );
  or2 U2211 ( .A1(n728), .A2(n729), .Z(n727) );
  and2 U2212 ( .A1(z2), .A2(n), .Z(n728) );
  or2 U2213 ( .A1(n730), .A2(n731), .Z(n729) );
  and2 U2214 ( .A1(i2), .A2(t), .Z(n730) );
  or2 U2215 ( .A1(n732), .A2(n733), .Z(n726) );
  and2 U2216 ( .A1(m), .A2(d3), .Z(n732) );
  or2 U2217 ( .A1(n734), .A2(n735), .Z(n733) );
  and2 U2218 ( .A1(c1), .A2(v), .Z(n734) );
  or2 U2219 ( .A1(n634), .A2(n635), .Z(n630) );
  and2 U2220 ( .A1(v1), .A2(q), .Z(n634) );
  or2 U2221 ( .A1(n636), .A2(n637), .Z(n635) );
  and2 U2222 ( .A1(o), .A2(r2), .Z(n636) );
  or2 U2223 ( .A1(n632), .A2(n633), .Z(n631) );
  and2 U2224 ( .A1(r), .A2(s1), .Z(n632) );
  and2 U2225 ( .A1(w), .A2(w0), .Z(n633) );
  or2 U2226 ( .A1(n640), .A2(n641), .Z(n639) );
  and2 U2227 ( .A1(n), .A2(y2), .Z(n640) );
  or2 U2228 ( .A1(n642), .A2(n643), .Z(n641) );
  and2 U2229 ( .A1(h2), .A2(t), .Z(n642) );
  or2 U2230 ( .A1(n644), .A2(n645), .Z(n638) );
  and2 U2231 ( .A1(m), .A2(c3), .Z(n644) );
  or2 U2232 ( .A1(n646), .A2(n647), .Z(n645) );
  and2 U2233 ( .A1(b1), .A2(v), .Z(n646) );
  or2 U2234 ( .A1(n581), .A2(n582), .Z(n577) );
  and2 U2235 ( .A1(p), .A2(p1), .Z(n581) );
  or2 U2236 ( .A1(n583), .A2(n584), .Z(n582) );
  and2 U2237 ( .A1(x2), .A2(n), .Z(n583) );
  or2 U2238 ( .A1(n579), .A2(n580), .Z(n578) );
  and2 U2239 ( .A1(q), .A2(r1), .Z(n579) );
  and2 U2240 ( .A1(w), .A2(v0), .Z(n580) );
  or2 U2241 ( .A1(n587), .A2(n588), .Z(n586) );
  and2 U2242 ( .A1(r), .A2(m1), .Z(n587) );
  or2 U2243 ( .A1(n589), .A2(n590), .Z(n588) );
  and2 U2244 ( .A1(f2), .A2(t), .Z(n589) );
  or2 U2245 ( .A1(n591), .A2(n592), .Z(n585) );
  and2 U2246 ( .A1(b3), .A2(m), .Z(n591) );
  or2 U2247 ( .A1(n593), .A2(n594), .Z(n592) );
  and2 U2248 ( .A1(a1), .A2(v), .Z(n593) );
  and2 U2249 ( .A1(z0), .A2(v), .Z(n503) );
  and2 U2250 ( .A1(p), .A2(q1), .Z(n502) );
  and2 U2251 ( .A1(t), .A2(e2), .Z(n510) );
  and2 U2252 ( .A1(q), .A2(n514), .Z(n513) );
  or2 U2253 ( .A1(n515), .A2(n516), .Z(n508) );
  or2 U2254 ( .A1(n517), .A2(n518), .Z(n516) );
  and2 U2255 ( .A1(s), .A2(n521), .Z(n515) );
  and2 U2256 ( .A1(o), .A2(n520), .Z(n517) );
  or2 U2257 ( .A1(n504), .A2(n505), .Z(n500) );
  and2 U2258 ( .A1(r), .A2(n1), .Z(n504) );
  or2 U2259 ( .A1(n506), .A2(n507), .Z(n505) );
  and2 U2260 ( .A1(w), .A2(l1), .Z(n506) );
  or2 U2261 ( .A1(n429), .A2(n430), .Z(n425) );
  and2 U2262 ( .A1(q4), .A2(q0), .Z(n429) );
  or2 U2263 ( .A1(n431), .A2(n432), .Z(n430) );
  and2 U2264 ( .A1(z3), .A2(o0), .Z(n431) );
  or2 U2265 ( .A1(n427), .A2(n428), .Z(n426) );
  and2 U2266 ( .A1(z4), .A2(t0), .Z(n427) );
  and2 U2267 ( .A1(u4), .A2(u0), .Z(n428) );
  or2 U2268 ( .A1(n435), .A2(n436), .Z(n434) );
  and2 U2269 ( .A1(l4), .A2(r0), .Z(n435) );
  or2 U2270 ( .A1(n437), .A2(n438), .Z(n436) );
  and2 U2271 ( .A1(t3), .A2(k0), .Z(n437) );
  or2 U2272 ( .A1(n439), .A2(n440), .Z(n433) );
  and2 U2273 ( .A1(i4), .A2(s0), .Z(n439) );
  or2 U2274 ( .A1(n441), .A2(n442), .Z(n440) );
  and2 U2275 ( .A1(c4), .A2(n0), .Z(n441) );
  or2 U2276 ( .A1(n356), .A2(n357), .Z(n352) );
  and2 U2277 ( .A1(v3), .A2(p0), .Z(n356) );
  or2 U2278 ( .A1(n358), .A2(n359), .Z(n357) );
  and2 U2279 ( .A1(y3), .A2(o0), .Z(n358) );
  or2 U2280 ( .A1(n354), .A2(n355), .Z(n353) );
  and2 U2281 ( .A1(y4), .A2(t0), .Z(n354) );
  and2 U2282 ( .A1(t4), .A2(u0), .Z(n355) );
  or2 U2283 ( .A1(n362), .A2(n363), .Z(n361) );
  and2 U2284 ( .A1(o3), .A2(l0), .Z(n362) );
  or2 U2285 ( .A1(n364), .A2(n365), .Z(n363) );
  and2 U2286 ( .A1(k0), .A2(s3), .Z(n364) );
  or2 U2287 ( .A1(n366), .A2(n367), .Z(n360) );
  and2 U2288 ( .A1(m0), .A2(h3), .Z(n366) );
  or2 U2289 ( .A1(n368), .A2(n369), .Z(n367) );
  and2 U2290 ( .A1(b4), .A2(n0), .Z(n368) );
  or2 U2291 ( .A1(n294), .A2(n295), .Z(n290) );
  and2 U2292 ( .A1(u3), .A2(p0), .Z(n294) );
  or2 U2293 ( .A1(n296), .A2(n297), .Z(n295) );
  and2 U2294 ( .A1(q0), .A2(n4), .Z(n296) );
  or2 U2295 ( .A1(n292), .A2(n293), .Z(n291) );
  and2 U2296 ( .A1(u0), .A2(s4), .Z(n292) );
  and2 U2297 ( .A1(x4), .A2(t0), .Z(n293) );
  or2 U2298 ( .A1(n300), .A2(n301), .Z(n299) );
  and2 U2299 ( .A1(n3), .A2(l0), .Z(n300) );
  or2 U2300 ( .A1(n302), .A2(n303), .Z(n301) );
  and2 U2301 ( .A1(r0), .A2(j4), .Z(n302) );
  or2 U2302 ( .A1(n304), .A2(n305), .Z(n298) );
  and2 U2303 ( .A1(m0), .A2(g3), .Z(n304) );
  or2 U2304 ( .A1(n306), .A2(n307), .Z(n305) );
  and2 U2305 ( .A1(n0), .A2(a4), .Z(n306) );
  or2 U2306 ( .A1(n1674), .A2(n1675), .Z(n1670) );
  and2 U2307 ( .A1(o0), .A2(r5), .Z(n1674) );
  or2 U2308 ( .A1(n1676), .A2(n1677), .Z(n1675) );
  and2 U2309 ( .A1(p0), .A2(m5), .Z(n1676) );
  or2 U2310 ( .A1(n1672), .A2(n1673), .Z(n1671) );
  and2 U2311 ( .A1(u0), .A2(r4), .Z(n1672) );
  and2 U2312 ( .A1(w4), .A2(t0), .Z(n1673) );
  or2 U2313 ( .A1(n1680), .A2(n1681), .Z(n1679) );
  and2 U2314 ( .A1(m4), .A2(q0), .Z(n1680) );
  or2 U2315 ( .A1(n1682), .A2(n1683), .Z(n1681) );
  and2 U2316 ( .A1(k0), .A2(q3), .Z(n1682) );
  or2 U2317 ( .A1(n1684), .A2(n1685), .Z(n1678) );
  and2 U2318 ( .A1(h4), .A2(r0), .Z(n1684) );
  or2 U2319 ( .A1(n1686), .A2(n1687), .Z(n1685) );
  and2 U2320 ( .A1(d4), .A2(s0), .Z(n1686) );
  and2 U2321 ( .A1(v4), .A2(t0), .Z(n1513) );
  and2 U2322 ( .A1(p0), .A2(n5), .Z(n1512) );
  and2 U2323 ( .A1(g4), .A2(r0), .Z(n1520) );
  and2 U2324 ( .A1(o0), .A2(n859), .Z(n1523) );
  or2 U2325 ( .A1(n1524), .A2(n1525), .Z(n1518) );
  or2 U2326 ( .A1(n1526), .A2(n1527), .Z(n1525) );
  and2 U2327 ( .A1(n960), .A2(q0), .Z(n1524) );
  and2 U2328 ( .A1(n653), .A2(m0), .Z(n1527) );
  or2 U2329 ( .A1(n1514), .A2(n1515), .Z(n1510) );
  and2 U2330 ( .A1(n0), .A2(q5), .Z(n1514) );
  or2 U2331 ( .A1(n1516), .A2(n1517), .Z(n1515) );
  and2 U2332 ( .A1(l3), .A2(l0), .Z(n1516) );
  and2 U2333 ( .A1(r1), .A2(n1953), .Z(n1799) );
  inv1 U2334 ( .I(v0), .ZN(n1965) );
  and2 U2335 ( .A1(v0), .A2(n1849), .Z(n1851) );
  and2 U2336 ( .A1(v0), .A2(n1854), .Z(n1855) );
  inv1 U2337 ( .I(n1853), .ZN(n1802) );
  or2 U2338 ( .A1(n1853), .A2(n1964), .Z(n1860) );
  inv1 U2339 ( .I(n1860), .ZN(n1858) );
  or2 U2340 ( .A1(n1860), .A2(n1963), .Z(n1862) );
  inv1 U2341 ( .I(n1862), .ZN(n1863) );
  inv1 U2342 ( .I(n1866), .ZN(n1867) );
  inv1 U2343 ( .I(a1), .ZN(n1827) );
  inv1 U2344 ( .I(n1810), .ZN(n1951) );
  or2 U2345 ( .A1(b), .A2(n876), .Z(n1447) );
  and2 U2346 ( .A1(n1837), .A2(n1726), .Z(n1838) );
  and2 U2347 ( .A1(n952), .A2(n1754), .Z(n1836) );
  and2 U2348 ( .A1(h1), .A2(n918), .Z(n952) );
  inv1 U2349 ( .I(h1), .ZN(n1842) );
  and2 U2350 ( .A1(n1879), .A2(n1726), .Z(n1841) );
  and2 U2351 ( .A1(n915), .A2(n1754), .Z(n1839) );
  and2 U2352 ( .A1(i1), .A2(n918), .Z(n915) );
  or2 U2353 ( .A1(n878), .A2(n879), .Z(n877) );
  and2 U2354 ( .A1(n521), .A2(n479), .Z(n879) );
  and2 U2355 ( .A1(j1), .A2(n480), .Z(n878) );
  and2 U2356 ( .A1(n1), .A2(n1454), .Z(n876) );
  and2 U2357 ( .A1(n1962), .A2(n695), .Z(n1454) );
  or2 U2358 ( .A1(n1881), .A2(n1880), .Z(n1883) );
  and2 U2359 ( .A1(n520), .A2(n1879), .Z(n1881) );
  inv1 U2360 ( .I(n1953), .ZN(n1880) );
  or2 U2361 ( .A1(n1894), .A2(n1886), .Z(n1882) );
  or2 U2362 ( .A1(n621), .A2(n1895), .Z(n1896) );
  and2 U2363 ( .A1(n1953), .A2(n1886), .Z(n1888) );
  and2 U2364 ( .A1(m1), .A2(n1), .Z(n1887) );
  or2 U2365 ( .A1(n1848), .A2(n693), .Z(n621) );
  or2 U2366 ( .A1(n497), .A2(n495), .Z(n693) );
  and2 U2367 ( .A1(n519), .A2(n1953), .Z(n1848) );
  and2 U2368 ( .A1(n520), .A2(n1953), .Z(n1847) );
  and2 U2369 ( .A1(n695), .A2(n1657), .Z(n623) );
  or2 U2370 ( .A1(n1776), .A2(b), .Z(n1969) );
  and2 U2371 ( .A1(n1657), .A2(n1775), .Z(n1776) );
  inv1 U2372 ( .I(l1), .ZN(n1775) );
  or2 U2373 ( .A1(r1), .A2(p1), .Z(n496) );
  or2 U2374 ( .A1(n491), .A2(q1), .Z(n490) );
  and2 U2375 ( .A1(n492), .A2(n493), .Z(n491) );
  or2 U2376 ( .A1(n494), .A2(n345), .Z(n493) );
  or2 U2377 ( .A1(n347), .A2(r1), .Z(n492) );
  or2 U2378 ( .A1(n482), .A2(n483), .Z(n415) );
  or2 U2379 ( .A1(b), .A2(n484), .Z(n483) );
  or2 U2380 ( .A1(n485), .A2(n486), .Z(n482) );
  and2 U2381 ( .A1(p1), .A2(q1), .Z(n484) );
  or2 U2382 ( .A1(q1), .A2(p1), .Z(n422) );
  or2 U2383 ( .A1(n418), .A2(r1), .Z(n417) );
  and2 U2384 ( .A1(n419), .A2(n420), .Z(n418) );
  or2 U2385 ( .A1(n347), .A2(p1), .Z(n419) );
  or2 U2386 ( .A1(n421), .A2(n345), .Z(n420) );
  or2 U2387 ( .A1(n497), .A2(d), .Z(n348) );
  or2 U2388 ( .A1(r1), .A2(q1), .Z(n349) );
  or2 U2389 ( .A1(n341), .A2(p1), .Z(n340) );
  and2 U2390 ( .A1(n342), .A2(n343), .Z(n341) );
  or2 U2391 ( .A1(n347), .A2(q1), .Z(n342) );
  or2 U2392 ( .A1(n344), .A2(n345), .Z(n343) );
  inv1 U2393 ( .I(n415), .ZN(n338) );
  and2 U2394 ( .A1(n283), .A2(n284), .Z(n281) );
  or2 U2395 ( .A1(s1), .A2(n1994), .Z(n283) );
  or2 U2396 ( .A1(n1996), .A2(n286), .Z(n284) );
  inv1 U2397 ( .I(b), .ZN(n1754) );
  and2 U2398 ( .A1(n1754), .A2(n1193), .Z(n282) );
  and2 U2399 ( .A1(n1754), .A2(n1207), .Z(n280) );
  or2 U2400 ( .A1(n1656), .A2(n623), .Z(n1207) );
  and2 U2401 ( .A1(n1658), .A2(v0), .Z(n1656) );
  and2 U2402 ( .A1(n1603), .A2(n1969), .Z(n1658) );
  inv1 U2403 ( .I(n1207), .ZN(n1193) );
  inv1 U2404 ( .I(b2), .ZN(n1113) );
  inv1 U2405 ( .I(n1112), .ZN(n1111) );
  or2 U2406 ( .A1(n1113), .A2(c2), .Z(n1112) );
  inv1 U2407 ( .I(n1039), .ZN(n1062) );
  and2 U2408 ( .A1(n1034), .A2(n574), .Z(n1033) );
  and2 U2409 ( .A1(n1035), .A2(n946), .Z(n1034) );
  or2 U2410 ( .A1(e2), .A2(n1036), .Z(n1035) );
  or2 U2411 ( .A1(n995), .A2(n996), .Z(n994) );
  and2 U2412 ( .A1(n909), .A2(n947), .Z(n996) );
  and2 U2413 ( .A1(f2), .A2(n946), .Z(n995) );
  or2 U2414 ( .A1(n574), .A2(t1), .Z(n992) );
  inv1 U2415 ( .I(n974), .ZN(n973) );
  or2 U2416 ( .A1(n942), .A2(n943), .Z(n941) );
  and2 U2417 ( .A1(h2), .A2(n945), .Z(n942) );
  inv1 U2418 ( .I(n944), .ZN(n943) );
  or2 U2419 ( .A1(n945), .A2(h2), .Z(n944) );
  or2 U2420 ( .A1(n574), .A2(u1), .Z(n939) );
  and2 U2421 ( .A1(n905), .A2(n574), .Z(n904) );
  or2 U2422 ( .A1(n906), .A2(n907), .Z(n905) );
  and2 U2423 ( .A1(n839), .A2(n873), .Z(n907) );
  and2 U2424 ( .A1(i2), .A2(n872), .Z(n906) );
  or2 U2425 ( .A1(n566), .A2(n867), .Z(n866) );
  or2 U2426 ( .A1(n868), .A2(n869), .Z(n867) );
  and2 U2427 ( .A1(j2), .A2(n871), .Z(n868) );
  inv1 U2428 ( .I(n870), .ZN(n869) );
  or2 U2429 ( .A1(k2), .A2(n836), .Z(n835) );
  and2 U2430 ( .A1(n617), .A2(h2), .Z(n616) );
  and2 U2431 ( .A1(f2), .A2(n618), .Z(n617) );
  or2 U2432 ( .A1(n574), .A2(b), .Z(n618) );
  and2 U2433 ( .A1(j2), .A2(i2), .Z(n615) );
  and2 U2434 ( .A1(l2), .A2(k2), .Z(n620) );
  and2 U2435 ( .A1(o2), .A2(m2), .Z(n619) );
  inv1 U2436 ( .I(n566), .ZN(n574) );
  or2 U2437 ( .A1(n479), .A2(n480), .Z(n477) );
  or2 U2438 ( .A1(a), .A2(n477), .Z(n478) );
  and2 U2439 ( .A1(q2), .A2(n275), .Z(n334) );
  inv1 U2440 ( .I(n1495), .ZN(n1492) );
  or2 U2441 ( .A1(n1238), .A2(n514), .Z(n1495) );
  and2 U2442 ( .A1(n703), .A2(n1494), .Z(n1493) );
  inv1 U2443 ( .I(z2), .ZN(n1494) );
  or2 U2444 ( .A1(n1895), .A2(b), .Z(n514) );
  and2 U2445 ( .A1(w2), .A2(n261), .Z(n1429) );
  inv1 U2446 ( .I(y2), .ZN(n703) );
  inv1 U2447 ( .I(n514), .ZN(n261) );
  and2 U2448 ( .A1(f3), .A2(n259), .Z(n968) );
  or2 U2449 ( .A1(n1952), .A2(z), .Z(n859) );
  inv1 U2450 ( .I(n863), .ZN(n860) );
  or2 U2451 ( .A1(n560), .A2(n859), .Z(n863) );
  and2 U2452 ( .A1(n557), .A2(n862), .Z(n861) );
  inv1 U2453 ( .I(o3), .ZN(n862) );
  and2 U2454 ( .A1(n3), .A2(n247), .Z(n830) );
  inv1 U2455 ( .I(l3), .ZN(n673) );
  inv1 U2456 ( .I(n3), .ZN(n557) );
  inv1 U2457 ( .I(n859), .ZN(n247) );
  and2 U2458 ( .A1(n1471), .A2(n1472), .Z(n1466) );
  or2 U2459 ( .A1(u3), .A2(n1473), .Z(n1471) );
  or2 U2460 ( .A1(n1167), .A2(n1425), .Z(n1472) );
  or2 U2461 ( .A1(n1368), .A2(n1369), .Z(n1367) );
  inv1 U2462 ( .I(n1370), .ZN(n1369) );
  and2 U2463 ( .A1(x3), .A2(n1322), .Z(n1319) );
  inv1 U2464 ( .I(n1322), .ZN(n1321) );
  and2 U2465 ( .A1(a4), .A2(n1164), .Z(n1161) );
  inv1 U2466 ( .I(n1164), .ZN(n1163) );
  and2 U2467 ( .A1(n1756), .A2(n1079), .Z(n1159) );
  and2 U2468 ( .A1(n1756), .A2(n1093), .Z(n1158) );
  or2 U2469 ( .A1(n1467), .A2(n650), .Z(n1093) );
  and2 U2470 ( .A1(n1469), .A2(n1470), .Z(n1467) );
  and2 U2471 ( .A1(r4), .A2(n1966), .Z(n1469) );
  inv1 U2472 ( .I(n1093), .ZN(n1079) );
  inv1 U2473 ( .I(e4), .ZN(n1015) );
  inv1 U2474 ( .I(d4), .ZN(n1016) );
  and2 U2475 ( .A1(d4), .A2(e4), .Z(n987) );
  inv1 U2476 ( .I(n986), .ZN(n985) );
  and2 U2477 ( .A1(n957), .A2(n394), .Z(n956) );
  and2 U2478 ( .A1(n958), .A2(n855), .Z(n957) );
  or2 U2479 ( .A1(g4), .A2(n959), .Z(n958) );
  or2 U2480 ( .A1(n923), .A2(n924), .Z(n922) );
  and2 U2481 ( .A1(n827), .A2(n856), .Z(n924) );
  and2 U2482 ( .A1(h4), .A2(n855), .Z(n923) );
  or2 U2483 ( .A1(n394), .A2(v3), .Z(n920) );
  inv1 U2484 ( .I(n888), .ZN(n887) );
  or2 U2485 ( .A1(n851), .A2(n852), .Z(n850) );
  and2 U2486 ( .A1(j4), .A2(n854), .Z(n851) );
  inv1 U2487 ( .I(n853), .ZN(n852) );
  or2 U2488 ( .A1(n854), .A2(j4), .Z(n853) );
  or2 U2489 ( .A1(n394), .A2(w3), .Z(n848) );
  and2 U2490 ( .A1(n823), .A2(n394), .Z(n822) );
  or2 U2491 ( .A1(n824), .A2(n825), .Z(n823) );
  and2 U2492 ( .A1(n664), .A2(n769), .Z(n825) );
  and2 U2493 ( .A1(k4), .A2(n770), .Z(n824) );
  or2 U2494 ( .A1(n386), .A2(n764), .Z(n763) );
  or2 U2495 ( .A1(n765), .A2(n766), .Z(n764) );
  and2 U2496 ( .A1(l4), .A2(n768), .Z(n765) );
  inv1 U2497 ( .I(n767), .ZN(n766) );
  or2 U2498 ( .A1(m4), .A2(n661), .Z(n660) );
  and2 U2499 ( .A1(n456), .A2(n4), .Z(n455) );
  and2 U2500 ( .A1(j4), .A2(n457), .Z(n456) );
  or2 U2501 ( .A1(n394), .A2(z), .Z(n457) );
  and2 U2502 ( .A1(o4), .A2(k4), .Z(n454) );
  and2 U2503 ( .A1(l4), .A2(h4), .Z(n459) );
  and2 U2504 ( .A1(q4), .A2(m4), .Z(n458) );
  or2 U2505 ( .A1(n960), .A2(n961), .Z(n386) );
  inv1 U2506 ( .I(n386), .ZN(n394) );
  and2 U2507 ( .A1(n1960), .A2(n1906), .Z(n1902) );
  and2 U2508 ( .A1(r4), .A2(n1906), .Z(n1907) );
  inv1 U2509 ( .I(n1905), .ZN(n1768) );
  inv1 U2510 ( .I(n1912), .ZN(n1910) );
  inv1 U2511 ( .I(n1914), .ZN(n1915) );
  inv1 U2512 ( .I(n1918), .ZN(n1919) );
  inv1 U2513 ( .I(w4), .ZN(n1813) );
  inv1 U2514 ( .I(n1774), .ZN(n1954) );
  and2 U2515 ( .A1(n1823), .A2(n1728), .Z(n1824) );
  and2 U2516 ( .A1(n1047), .A2(d5), .Z(n1822) );
  inv1 U2517 ( .I(d5), .ZN(n1835) );
  and2 U2518 ( .A1(n1936), .A2(n1728), .Z(n1834) );
  and2 U2519 ( .A1(n1047), .A2(e5), .Z(n1832) );
  or2 U2520 ( .A1(f5), .A2(g5), .Z(n1003) );
  and2 U2521 ( .A1(f5), .A2(n981), .Z(n999) );
  or2 U2522 ( .A1(n747), .A2(n1699), .Z(n1011) );
  or2 U2523 ( .A1(m5), .A2(n746), .Z(n1699) );
  or2 U2524 ( .A1(n746), .A2(n1468), .Z(n1010) );
  or2 U2525 ( .A1(n5), .A2(m5), .Z(n1468) );
  or2 U2526 ( .A1(n961), .A2(n650), .Z(n977) );
  and2 U2527 ( .A1(f5), .A2(n982), .Z(n979) );
  inv1 U2528 ( .I(j5), .ZN(n883) );
  inv1 U2529 ( .I(k5), .ZN(n846) );
  or2 U2530 ( .A1(n844), .A2(k5), .Z(n843) );
  and2 U2531 ( .A1(n884), .A2(n1756), .Z(n841) );
  or2 U2532 ( .A1(n846), .A2(j5), .Z(n884) );
  inv1 U2533 ( .I(n1945), .ZN(n1952) );
  or2 U2534 ( .A1(n1791), .A2(n1790), .Z(n1945) );
  or2 U2535 ( .A1(l5), .A2(n5), .Z(n1791) );
  or2 U2536 ( .A1(n1956), .A2(z), .Z(n1790) );
  and2 U2537 ( .A1(n1749), .A2(n1932), .Z(n1933) );
  or2 U2538 ( .A1(n1931), .A2(n1843), .Z(n1932) );
  inv1 U2539 ( .I(n1937), .ZN(n1939) );
  and2 U2540 ( .A1(m5), .A2(n5), .Z(n1938) );
  inv1 U2541 ( .I(z), .ZN(n1756) );
  or2 U2542 ( .A1(n1846), .A2(n742), .Z(n648) );
  or2 U2543 ( .A1(n538), .A2(n536), .Z(n742) );
  or2 U2544 ( .A1(n1844), .A2(n1931), .Z(n1845) );
  inv1 U2545 ( .I(n1010), .ZN(n650) );
  and2 U2546 ( .A1(n1696), .A2(n1957), .Z(n1770) );
  and2 U2547 ( .A1(n1956), .A2(n747), .Z(n1696) );
  or2 U2548 ( .A1(r5), .A2(p5), .Z(n537) );
  or2 U2549 ( .A1(n532), .A2(q5), .Z(n531) );
  and2 U2550 ( .A1(n533), .A2(n534), .Z(n532) );
  or2 U2551 ( .A1(n535), .A2(n378), .Z(n534) );
  or2 U2552 ( .A1(n380), .A2(r5), .Z(n533) );
  or2 U2553 ( .A1(n523), .A2(n524), .Z(n444) );
  or2 U2554 ( .A1(z), .A2(n525), .Z(n524) );
  or2 U2555 ( .A1(n526), .A2(n527), .Z(n523) );
  and2 U2556 ( .A1(p5), .A2(q5), .Z(n525) );
  or2 U2557 ( .A1(q5), .A2(p5), .Z(n451) );
  or2 U2558 ( .A1(n447), .A2(r5), .Z(n446) );
  and2 U2559 ( .A1(n448), .A2(n449), .Z(n447) );
  or2 U2560 ( .A1(n380), .A2(p5), .Z(n448) );
  or2 U2561 ( .A1(n450), .A2(n378), .Z(n449) );
  or2 U2562 ( .A1(n538), .A2(b0), .Z(n381) );
  or2 U2563 ( .A1(r5), .A2(q5), .Z(n382) );
  or2 U2564 ( .A1(n374), .A2(p5), .Z(n373) );
  and2 U2565 ( .A1(n375), .A2(n376), .Z(n374) );
  or2 U2566 ( .A1(n380), .A2(q5), .Z(n375) );
  or2 U2567 ( .A1(n377), .A2(n378), .Z(n376) );
  inv1 U2568 ( .I(n444), .ZN(n371) );
  inv1 U2569 ( .I(n1653), .ZN(n1652) );
  or2 U2570 ( .A1(n1654), .A2(n1655), .Z(n1653) );
  or2 U2571 ( .A1(b1), .A2(c1), .Z(n1655) );
  and2 U2572 ( .A1(n1440), .A2(n1297), .Z(n1300) );
  or2 U2573 ( .A1(n1441), .A2(s1), .Z(n1440) );
  or2 U2574 ( .A1(t1), .A2(u1), .Z(n1441) );
  or2 U2575 ( .A1(v1), .A2(n1300), .Z(n1299) );
  or2 U2576 ( .A1(x1), .A2(w1), .Z(n1298) );
  and2 U2577 ( .A1(n1325), .A2(n1170), .Z(n1173) );
  or2 U2578 ( .A1(n1326), .A2(u3), .Z(n1325) );
  or2 U2579 ( .A1(v3), .A2(w3), .Z(n1326) );
  or2 U2580 ( .A1(x3), .A2(n1173), .Z(n1172) );
  or2 U2581 ( .A1(z3), .A2(y3), .Z(n1171) );
  or2 U2582 ( .A1(a3), .A2(n705), .Z(n704) );
  or2 U2583 ( .A1(z2), .A2(e3), .Z(n706) );
  inv1 U2584 ( .I(n348), .ZN(n346) );
  and2 U2585 ( .A1(n1648), .A2(n1969), .Z(n1647) );
  or2 U2586 ( .A1(n1649), .A2(p1), .Z(n1648) );
  or2 U2587 ( .A1(n1652), .A2(q1), .Z(n1650) );
  and2 U2588 ( .A1(n1964), .A2(n1963), .Z(n1646) );
  or2 U2589 ( .A1(b1), .A2(a1), .Z(n1665) );
  or2 U2590 ( .A1(d1), .A2(c1), .Z(n1664) );
  or2 U2591 ( .A1(x0), .A2(w0), .Z(n1667) );
  or2 U2592 ( .A1(z0), .A2(y0), .Z(n1666) );
  and2 U2593 ( .A1(n1482), .A2(n1966), .Z(n1481) );
  or2 U2594 ( .A1(n1483), .A2(p5), .Z(n1482) );
  and2 U2595 ( .A1(n1484), .A2(n1811), .Z(n1483) );
  and2 U2596 ( .A1(n1959), .A2(n1958), .Z(n1477) );
  or2 U2597 ( .A1(t4), .A2(s4), .Z(n1574) );
  or2 U2598 ( .A1(v4), .A2(u4), .Z(n1573) );
  or2 U2599 ( .A1(x4), .A2(w4), .Z(n1576) );
  or2 U2600 ( .A1(z4), .A2(y4), .Z(n1575) );
  or2 U2601 ( .A1(o3), .A2(n557), .Z(n1535) );
  or2 U2602 ( .A1(t3), .A2(q3), .Z(n1536) );
  or2 U2603 ( .A1(r3), .A2(s3), .Z(n1534) );
  inv1 U2604 ( .I(n381), .ZN(n379) );
  and2 U2605 ( .A1(o2), .A2(s), .Z(n804) );
  and2 U2606 ( .A1(u), .A2(g2), .Z(n810) );
  and2 U2607 ( .A1(a3), .A2(n), .Z(n814) );
  and2 U2608 ( .A1(z1), .A2(p), .Z(n725) );
  and2 U2609 ( .A1(m2), .A2(s), .Z(n731) );
  and2 U2610 ( .A1(u), .A2(d2), .Z(n735) );
  and2 U2611 ( .A1(y1), .A2(p), .Z(n637) );
  and2 U2612 ( .A1(l2), .A2(s), .Z(n643) );
  and2 U2613 ( .A1(u), .A2(c2), .Z(n647) );
  and2 U2614 ( .A1(o), .A2(q2), .Z(n584) );
  and2 U2615 ( .A1(k2), .A2(s), .Z(n590) );
  and2 U2616 ( .A1(u), .A2(b2), .Z(n594) );
  and2 U2617 ( .A1(m), .A2(n519), .Z(n518) );
  and2 U2618 ( .A1(n), .A2(w2), .Z(n507) );
  and2 U2619 ( .A1(w3), .A2(p0), .Z(n432) );
  and2 U2620 ( .A1(l0), .A2(p3), .Z(n438) );
  and2 U2621 ( .A1(m0), .A2(i3), .Z(n442) );
  and2 U2622 ( .A1(o4), .A2(q0), .Z(n359) );
  and2 U2623 ( .A1(k4), .A2(r0), .Z(n365) );
  and2 U2624 ( .A1(f4), .A2(s0), .Z(n369) );
  and2 U2625 ( .A1(x3), .A2(o0), .Z(n297) );
  and2 U2626 ( .A1(k0), .A2(r3), .Z(n303) );
  and2 U2627 ( .A1(s0), .A2(e4), .Z(n307) );
  and2 U2628 ( .A1(n0), .A2(p5), .Z(n1677) );
  and2 U2629 ( .A1(m3), .A2(l0), .Z(n1683) );
  and2 U2630 ( .A1(m0), .A2(f3), .Z(n1687) );
  and2 U2631 ( .A1(n1528), .A2(n1529), .Z(n653) );
  and2 U2632 ( .A1(s3), .A2(t3), .Z(n1529) );
  and2 U2633 ( .A1(r3), .A2(n1530), .Z(n1528) );
  and2 U2634 ( .A1(p3), .A2(q3), .Z(n1530) );
  and2 U2635 ( .A1(n751), .A2(k0), .Z(n1526) );
  and2 U2636 ( .A1(u0), .A2(l5), .Z(n1517) );
  inv1 U2637 ( .I(z0), .ZN(n1825) );
  and2 U2638 ( .A1(n1969), .A2(n1805), .Z(n1808) );
  inv1 U2639 ( .I(n2036), .ZN(n1805) );
  and2 U2640 ( .A1(n1953), .A2(n1806), .Z(n1807) );
  and2 U2641 ( .A1(v0), .A2(r1), .Z(n1806) );
  inv1 U2642 ( .I(n876), .ZN(n918) );
  inv1 U2643 ( .I(m1), .ZN(n1962) );
  and2 U2644 ( .A1(n1), .A2(n694), .Z(n495) );
  and2 U2645 ( .A1(m1), .A2(n695), .Z(n694) );
  inv1 U2646 ( .I(n700), .ZN(n519) );
  or2 U2647 ( .A1(n701), .A2(n702), .Z(n700) );
  or2 U2648 ( .A1(b3), .A2(n706), .Z(n701) );
  or2 U2649 ( .A1(n703), .A2(n704), .Z(n702) );
  and2 U2650 ( .A1(n346), .A2(p1), .Z(n494) );
  and2 U2651 ( .A1(n487), .A2(n1961), .Z(n486) );
  inv1 U2652 ( .I(n422), .ZN(n487) );
  and2 U2653 ( .A1(r1), .A2(n422), .Z(n485) );
  and2 U2654 ( .A1(n346), .A2(q1), .Z(n421) );
  or2 U2655 ( .A1(n495), .A2(e), .Z(n345) );
  and2 U2656 ( .A1(n346), .A2(r1), .Z(n344) );
  inv1 U2657 ( .I(n345), .ZN(n347) );
  or2 U2658 ( .A1(n1996), .A2(n1633), .Z(n1632) );
  or2 U2659 ( .A1(n1818), .A2(s1), .Z(n1634) );
  and2 U2660 ( .A1(n1796), .A2(n1985), .Z(n1503) );
  inv1 U2661 ( .I(n1444), .ZN(n1796) );
  and2 U2662 ( .A1(n1402), .A2(n1985), .Z(n1438) );
  and2 U2663 ( .A1(n1357), .A2(n1818), .Z(n1399) );
  inv1 U2664 ( .I(x1), .ZN(n1303) );
  or2 U2665 ( .A1(n1354), .A2(n1355), .Z(n1353) );
  and2 U2666 ( .A1(n1302), .A2(n1818), .Z(n1354) );
  and2 U2667 ( .A1(n1251), .A2(n1985), .Z(n1293) );
  and2 U2668 ( .A1(n1206), .A2(n1985), .Z(n1248) );
  or2 U2669 ( .A1(n1200), .A2(n1201), .Z(n1199) );
  or2 U2670 ( .A1(p1), .A2(l), .Z(n1037) );
  inv1 U2671 ( .I(f2), .ZN(n947) );
  inv1 U2672 ( .I(n909), .ZN(n946) );
  or2 U2673 ( .A1(n946), .A2(n947), .Z(n945) );
  inv1 U2674 ( .I(n839), .ZN(n872) );
  inv1 U2675 ( .I(i2), .ZN(n873) );
  or2 U2676 ( .A1(n871), .A2(j2), .Z(n870) );
  or2 U2677 ( .A1(n872), .A2(n873), .Z(n871) );
  inv1 U2678 ( .I(n686), .ZN(n788) );
  inv1 U2679 ( .I(m2), .ZN(n573) );
  and2 U2680 ( .A1(n1603), .A2(n1965), .Z(n1789) );
  inv1 U2681 ( .I(x2), .ZN(n1284) );
  inv1 U2682 ( .I(c3), .ZN(n1058) );
  inv1 U2683 ( .I(d3), .ZN(n1029) );
  or2 U2684 ( .A1(c3), .A2(d3), .Z(n705) );
  or2 U2685 ( .A1(r4), .A2(n1955), .Z(n1578) );
  and2 U2686 ( .A1(n1470), .A2(n1960), .Z(n1795) );
  inv1 U2687 ( .I(n472), .ZN(n672) );
  inv1 U2688 ( .I(m3), .ZN(n612) );
  or2 U2689 ( .A1(l3), .A2(m3), .Z(n560) );
  inv1 U2690 ( .I(j3), .ZN(n470) );
  inv1 U2691 ( .I(k3), .ZN(n474) );
  inv1 U2692 ( .I(r3), .ZN(n325) );
  inv1 U2693 ( .I(s3), .ZN(n252) );
  inv1 U2694 ( .I(u3), .ZN(n1425) );
  and2 U2695 ( .A1(n1798), .A2(n1820), .Z(n1372) );
  inv1 U2696 ( .I(n1329), .ZN(n1798) );
  and2 U2697 ( .A1(n1274), .A2(n1820), .Z(n1323) );
  and2 U2698 ( .A1(n1225), .A2(n1820), .Z(n1271) );
  inv1 U2699 ( .I(z3), .ZN(n1176) );
  and2 U2700 ( .A1(n1175), .A2(n1820), .Z(n1222) );
  and2 U2701 ( .A1(n1128), .A2(n1820), .Z(n1165) );
  and2 U2702 ( .A1(n1092), .A2(n1820), .Z(n1125) );
  inv1 U2703 ( .I(n1570), .ZN(n1470) );
  or2 U2704 ( .A1(n1571), .A2(n1572), .Z(n1570) );
  or2 U2705 ( .A1(n1575), .A2(n1576), .Z(n1571) );
  or2 U2706 ( .A1(n1573), .A2(n1574), .Z(n1572) );
  and2 U2707 ( .A1(n1089), .A2(n1820), .Z(n1086) );
  or2 U2708 ( .A1(p5), .A2(j0), .Z(n1537) );
  inv1 U2709 ( .I(h4), .ZN(n856) );
  inv1 U2710 ( .I(n827), .ZN(n855) );
  or2 U2711 ( .A1(n855), .A2(n856), .Z(n854) );
  inv1 U2712 ( .I(n664), .ZN(n770) );
  inv1 U2713 ( .I(k4), .ZN(n769) );
  or2 U2714 ( .A1(n768), .A2(l4), .Z(n767) );
  or2 U2715 ( .A1(n769), .A2(n770), .Z(n768) );
  inv1 U2716 ( .I(n546), .ZN(n602) );
  inv1 U2717 ( .I(o4), .ZN(n392) );
  inv1 U2718 ( .I(v4), .ZN(n1811) );
  or2 U2719 ( .A1(n1924), .A2(n1814), .Z(n1815) );
  inv1 U2720 ( .I(y4), .ZN(n1814) );
  and2 U2721 ( .A1(n1966), .A2(n1771), .Z(n1772) );
  inv1 U2722 ( .I(n2012), .ZN(n1771) );
  and2 U2723 ( .A1(n1698), .A2(r5), .Z(n1692) );
  inv1 U2724 ( .I(n743), .ZN(n536) );
  or2 U2725 ( .A1(n1956), .A2(n745), .Z(n743) );
  or2 U2726 ( .A1(n746), .A2(n747), .Z(n745) );
  inv1 U2727 ( .I(n1531), .ZN(n751) );
  or2 U2728 ( .A1(n1532), .A2(n1533), .Z(n1531) );
  or2 U2729 ( .A1(p3), .A2(n1536), .Z(n1532) );
  or2 U2730 ( .A1(n1534), .A2(n1535), .Z(n1533) );
  inv1 U2731 ( .I(n653), .ZN(n1843) );
  inv1 U2732 ( .I(m5), .ZN(n1956) );
  and2 U2733 ( .A1(n379), .A2(p5), .Z(n535) );
  and2 U2734 ( .A1(n528), .A2(n1955), .Z(n527) );
  inv1 U2735 ( .I(n451), .ZN(n528) );
  and2 U2736 ( .A1(r5), .A2(n451), .Z(n526) );
  and2 U2737 ( .A1(n379), .A2(q5), .Z(n450) );
  and2 U2738 ( .A1(n379), .A2(r5), .Z(n377) );
  or2 U2739 ( .A1(n536), .A2(c0), .Z(n378) );
  inv1 U2740 ( .I(n378), .ZN(n380) );
  inv1 U2741 ( .I(d1), .ZN(n1068) );
  or2 U2742 ( .A1(n785), .A2(n786), .Z(n784) );
  and2 U2743 ( .A1(n686), .A2(n787), .Z(n786) );
  and2 U2744 ( .A1(l2), .A2(n788), .Z(n785) );
  inv1 U2745 ( .I(l2), .ZN(n787) );
  and2 U2746 ( .A1(n276), .A2(n2023), .Z(n267) );
  and2 U2747 ( .A1(n271), .A2(n272), .Z(n270) );
  or2 U2748 ( .A1(n1390), .A2(n1978), .Z(n1609) );
  or2 U2749 ( .A1(n1384), .A2(n1338), .Z(n1383) );
  and2 U2750 ( .A1(n1385), .A2(n1978), .Z(n1384) );
  inv1 U2751 ( .I(n1151), .ZN(n1385) );
  and2 U2752 ( .A1(n1337), .A2(n1338), .Z(n1336) );
  or2 U2753 ( .A1(n1342), .A2(n1343), .Z(n1340) );
  and2 U2754 ( .A1(n1978), .A2(n1285), .Z(n1342) );
  and2 U2755 ( .A1(w2), .A2(n2023), .Z(n1343) );
  inv1 U2756 ( .I(n1148), .ZN(n1142) );
  and2 U2757 ( .A1(n1139), .A2(n2023), .Z(n1135) );
  and2 U2758 ( .A1(n514), .A2(n1978), .Z(n1018) );
  and2 U2759 ( .A1(n937), .A2(n2038), .Z(n930) );
  and2 U2760 ( .A1(n933), .A2(n934), .Z(n932) );
  or2 U2761 ( .A1(n901), .A2(n259), .Z(n897) );
  and2 U2762 ( .A1(n473), .A2(n259), .Z(n779) );
  or2 U2763 ( .A1(n677), .A2(n678), .Z(n675) );
  and2 U2764 ( .A1(n1971), .A2(n611), .Z(n677) );
  and2 U2765 ( .A1(l3), .A2(n2037), .Z(n678) );
  or2 U2766 ( .A1(n2037), .A2(q3), .Z(n409) );
  and2 U2767 ( .A1(n859), .A2(n1971), .Z(n246) );
  or2 U2768 ( .A1(n1418), .A2(n1419), .Z(n1417) );
  and2 U2769 ( .A1(v3), .A2(n1421), .Z(n1418) );
  inv1 U2770 ( .I(n1420), .ZN(n1419) );
  or2 U2771 ( .A1(n599), .A2(n600), .Z(n598) );
  and2 U2772 ( .A1(n546), .A2(n601), .Z(n600) );
  and2 U2773 ( .A1(n4), .A2(n602), .Z(n599) );
  inv1 U2774 ( .I(n4), .ZN(n601) );
  inv1 U2775 ( .I(z4), .ZN(n1261) );
  or2 U2776 ( .A1(n1005), .A2(n977), .Z(n1967) );
  and2 U2777 ( .A1(h5), .A2(n1009), .Z(n1007) );
  or2 U2778 ( .A1(n805), .A2(n806), .Z(n795) );
  or2 U2779 ( .A1(n797), .A2(n798), .Z(n796) );
  or2 U2780 ( .A1(n726), .A2(n727), .Z(n716) );
  or2 U2781 ( .A1(n718), .A2(n719), .Z(n717) );
  or2 U2782 ( .A1(n638), .A2(n639), .Z(n628) );
  or2 U2783 ( .A1(n630), .A2(n631), .Z(n629) );
  or2 U2784 ( .A1(n585), .A2(n586), .Z(n575) );
  or2 U2785 ( .A1(n577), .A2(n578), .Z(n576) );
  or2 U2786 ( .A1(n500), .A2(n501), .Z(n499) );
  or2 U2787 ( .A1(n502), .A2(n503), .Z(n501) );
  or2 U2788 ( .A1(n433), .A2(n434), .Z(n423) );
  or2 U2789 ( .A1(n425), .A2(n426), .Z(n424) );
  or2 U2790 ( .A1(n360), .A2(n361), .Z(n350) );
  or2 U2791 ( .A1(n352), .A2(n353), .Z(n351) );
  or2 U2792 ( .A1(n298), .A2(n299), .Z(n288) );
  or2 U2793 ( .A1(n290), .A2(n291), .Z(n289) );
  or2 U2794 ( .A1(n1678), .A2(n1679), .Z(n1668) );
  or2 U2795 ( .A1(n1670), .A2(n1671), .Z(n1669) );
  or2 U2796 ( .A1(n1510), .A2(n1511), .Z(n1509) );
  or2 U2797 ( .A1(n1512), .A2(n1513), .Z(n1511) );
  or2 U2798 ( .A1(n1851), .A2(n1850), .Z(n1852) );
  and2 U2799 ( .A1(n1965), .A2(n1854), .Z(n1850) );
  or2 U2800 ( .A1(n1855), .A2(w0), .Z(n1856) );
  and2 U2801 ( .A1(n1853), .A2(n1951), .Z(n1857) );
  and2 U2802 ( .A1(n1860), .A2(n1803), .Z(n1358) );
  or2 U2803 ( .A1(n1802), .A2(x0), .Z(n1803) );
  and2 U2804 ( .A1(n1951), .A2(n1859), .Z(n1861) );
  and2 U2805 ( .A1(n1951), .A2(n1866), .Z(n1865) );
  or2 U2806 ( .A1(n1863), .A2(z0), .Z(n1864) );
  or2 U2807 ( .A1(n1867), .A2(a1), .Z(n1868) );
  and2 U2808 ( .A1(n1951), .A2(n1873), .Z(n1869) );
  and2 U2809 ( .A1(n1874), .A2(n1875), .Z(i6) );
  or2 U2810 ( .A1(n1870), .A2(b1), .Z(n1871) );
  and2 U2811 ( .A1(n1878), .A2(n1877), .Z(j6) );
  or2 U2812 ( .A1(n1876), .A2(c1), .Z(n1877) );
  and2 U2813 ( .A1(n1886), .A2(n1836), .Z(n948) );
  and2 U2814 ( .A1(n1842), .A2(n1838), .Z(n949) );
  and2 U2815 ( .A1(n2028), .A2(n1839), .Z(n910) );
  and2 U2816 ( .A1(n1842), .A2(n1841), .Z(n911) );
  or2 U2817 ( .A1(n623), .A2(n876), .Z(n875) );
  and2 U2818 ( .A1(n877), .A2(n1754), .Z(n874) );
  inv1 U2819 ( .I(n1884), .ZN(n1885) );
  and2 U2820 ( .A1(n1883), .A2(n1882), .Z(n1884) );
  or2 U2821 ( .A1(n1888), .A2(n1887), .Z(n1899) );
  or2 U2822 ( .A1(n623), .A2(n624), .Z(n622) );
  and2 U2823 ( .A1(n1879), .A2(n1847), .Z(n624) );
  and2 U2824 ( .A1(n489), .A2(n490), .Z(n481) );
  or2 U2825 ( .A1(n348), .A2(n496), .Z(n489) );
  and2 U2826 ( .A1(n416), .A2(n417), .Z(n414) );
  or2 U2827 ( .A1(n348), .A2(n422), .Z(n416) );
  and2 U2828 ( .A1(n339), .A2(n340), .Z(n337) );
  or2 U2829 ( .A1(n348), .A2(n349), .Z(n339) );
  and2 U2830 ( .A1(w2), .A2(n280), .Z(n279) );
  and2 U2831 ( .A1(n281), .A2(n282), .Z(n278) );
  and2 U2832 ( .A1(n1625), .A2(n1626), .Z(a7) );
  or2 U2833 ( .A1(n1193), .A2(x2), .Z(n1626) );
  and2 U2834 ( .A1(y2), .A2(n280), .Z(n1497) );
  or2 U2835 ( .A1(n1430), .A2(n1431), .Z(c7) );
  and2 U2836 ( .A1(z2), .A2(n1207), .Z(n1430) );
  and2 U2837 ( .A1(a3), .A2(n1207), .Z(n1391) );
  and2 U2838 ( .A1(b3), .A2(n1207), .Z(n1344) );
  and2 U2839 ( .A1(c3), .A2(n280), .Z(n1287) );
  and2 U2840 ( .A1(d3), .A2(n1207), .Z(n1240) );
  and2 U2841 ( .A1(e3), .A2(n1207), .Z(n1189) );
  or2 U2842 ( .A1(n1110), .A2(n1111), .Z(n1109) );
  and2 U2843 ( .A1(c2), .A2(n1113), .Z(n1110) );
  and2 U2844 ( .A1(n1061), .A2(n1062), .Z(n1060) );
  or2 U2845 ( .A1(n1063), .A2(d2), .Z(n1061) );
  and2 U2846 ( .A1(s1), .A2(n566), .Z(n1031) );
  or2 U2847 ( .A1(b), .A2(n1033), .Z(n1032) );
  and2 U2848 ( .A1(n992), .A2(n993), .Z(n991) );
  or2 U2849 ( .A1(n566), .A2(n994), .Z(n993) );
  and2 U2850 ( .A1(n972), .A2(n973), .Z(n971) );
  or2 U2851 ( .A1(g2), .A2(n975), .Z(n972) );
  and2 U2852 ( .A1(n939), .A2(n940), .Z(n938) );
  or2 U2853 ( .A1(n566), .A2(n941), .Z(n940) );
  and2 U2854 ( .A1(v1), .A2(n566), .Z(n902) );
  or2 U2855 ( .A1(b), .A2(n904), .Z(n903) );
  and2 U2856 ( .A1(n865), .A2(n866), .Z(n864) );
  or2 U2857 ( .A1(n574), .A2(w1), .Z(n865) );
  and2 U2858 ( .A1(x1), .A2(n566), .Z(n831) );
  or2 U2859 ( .A1(b), .A2(n833), .Z(n832) );
  or2 U2860 ( .A1(n574), .A2(z1), .Z(n680) );
  and2 U2861 ( .A1(n619), .A2(n620), .Z(n613) );
  and2 U2862 ( .A1(n615), .A2(n616), .Z(n614) );
  or2 U2863 ( .A1(n574), .A2(a2), .Z(n564) );
  inv1 U2864 ( .I(n478), .ZN(n475) );
  and2 U2865 ( .A1(p2), .A2(n477), .Z(n476) );
  and2 U2866 ( .A1(n411), .A2(n261), .Z(x7) );
  and2 U2867 ( .A1(n412), .A2(n413), .Z(n411) );
  or2 U2868 ( .A1(q2), .A2(n1979), .Z(n412) );
  or2 U2869 ( .A1(n330), .A2(r2), .Z(n329) );
  inv1 U2870 ( .I(n331), .ZN(n328) );
  and2 U2871 ( .A1(n1492), .A2(n1493), .Z(n1490) );
  and2 U2872 ( .A1(n2022), .A2(n514), .Z(n1491) );
  and2 U2873 ( .A1(z2), .A2(x2), .Z(n1427) );
  and2 U2874 ( .A1(n1429), .A2(y2), .Z(n1428) );
  and2 U2875 ( .A1(n988), .A2(n247), .Z(m8) );
  and2 U2876 ( .A1(n989), .A2(n990), .Z(n988) );
  or2 U2877 ( .A1(f3), .A2(n2048), .Z(n989) );
  and2 U2878 ( .A1(n962), .A2(n247), .Z(n8) );
  and2 U2879 ( .A1(n860), .A2(n861), .Z(n857) );
  and2 U2880 ( .A1(n2037), .A2(n859), .Z(n858) );
  and2 U2881 ( .A1(m3), .A2(l3), .Z(n828) );
  and2 U2882 ( .A1(n830), .A2(o3), .Z(n829) );
  and2 U2883 ( .A1(n1158), .A2(l3), .Z(n1465) );
  and2 U2884 ( .A1(n1466), .A2(n1159), .Z(n1464) );
  and2 U2885 ( .A1(n1158), .A2(n3), .Z(n1366) );
  and2 U2886 ( .A1(o3), .A2(n1093), .Z(n1315) );
  and2 U2887 ( .A1(p3), .A2(n1093), .Z(n1263) );
  and2 U2888 ( .A1(q3), .A2(n1093), .Z(n1212) );
  and2 U2889 ( .A1(n1158), .A2(r3), .Z(n1157) );
  and2 U2890 ( .A1(s3), .A2(n1093), .Z(n1117) );
  and2 U2891 ( .A1(t3), .A2(n1093), .Z(n1075) );
  or2 U2892 ( .A1(n1013), .A2(n1014), .Z(n1012) );
  and2 U2893 ( .A1(e4), .A2(n1016), .Z(n1013) );
  and2 U2894 ( .A1(d4), .A2(n1015), .Z(n1014) );
  and2 U2895 ( .A1(n984), .A2(n985), .Z(n983) );
  or2 U2896 ( .A1(n987), .A2(f4), .Z(n984) );
  and2 U2897 ( .A1(u3), .A2(n386), .Z(n954) );
  or2 U2898 ( .A1(z), .A2(n956), .Z(n955) );
  and2 U2899 ( .A1(n920), .A2(n921), .Z(n919) );
  or2 U2900 ( .A1(n386), .A2(n922), .Z(n921) );
  and2 U2901 ( .A1(n886), .A2(n887), .Z(n885) );
  or2 U2902 ( .A1(i4), .A2(n889), .Z(n886) );
  and2 U2903 ( .A1(n848), .A2(n849), .Z(n847) );
  or2 U2904 ( .A1(n386), .A2(n850), .Z(n849) );
  and2 U2905 ( .A1(x3), .A2(n386), .Z(n820) );
  or2 U2906 ( .A1(z), .A2(n822), .Z(n821) );
  and2 U2907 ( .A1(n762), .A2(n763), .Z(n761) );
  or2 U2908 ( .A1(n394), .A2(y3), .Z(n762) );
  and2 U2909 ( .A1(z3), .A2(n386), .Z(n656) );
  or2 U2910 ( .A1(z), .A2(n658), .Z(n657) );
  or2 U2911 ( .A1(n595), .A2(z), .Z(u9) );
  and2 U2912 ( .A1(n596), .A2(n597), .Z(n595) );
  or2 U2913 ( .A1(n394), .A2(a4), .Z(n596) );
  or2 U2914 ( .A1(n386), .A2(n598), .Z(n597) );
  or2 U2915 ( .A1(n394), .A2(b4), .Z(n540) );
  and2 U2916 ( .A1(n458), .A2(n459), .Z(n452) );
  and2 U2917 ( .A1(n454), .A2(n455), .Z(n453) );
  or2 U2918 ( .A1(n394), .A2(c4), .Z(n384) );
  or2 U2919 ( .A1(n1903), .A2(n1902), .Z(n1904) );
  and2 U2920 ( .A1(r4), .A2(n1901), .Z(n1903) );
  or2 U2921 ( .A1(n1907), .A2(s4), .Z(n1908) );
  and2 U2922 ( .A1(n1905), .A2(n1954), .Z(n1909) );
  and2 U2923 ( .A1(n1912), .A2(n1769), .Z(n1688) );
  or2 U2924 ( .A1(n1768), .A2(t4), .Z(n1769) );
  and2 U2925 ( .A1(n1954), .A2(n1911), .Z(n1913) );
  and2 U2926 ( .A1(n1954), .A2(n1918), .Z(n1917) );
  or2 U2927 ( .A1(n1915), .A2(v4), .Z(n1916) );
  or2 U2928 ( .A1(n1919), .A2(w4), .Z(n1920) );
  and2 U2929 ( .A1(n1954), .A2(n1925), .Z(n1921) );
  and2 U2930 ( .A1(n1926), .A2(n1927), .Z(e10) );
  or2 U2931 ( .A1(n1922), .A2(x4), .Z(n1923) );
  inv1 U2932 ( .I(n1925), .ZN(n1922) );
  and2 U2933 ( .A1(n1930), .A2(n1929), .Z(f10) );
  or2 U2934 ( .A1(n1928), .A2(y4), .Z(n1929) );
  and2 U2935 ( .A1(n1954), .A2(n1725), .Z(n1930) );
  inv1 U2936 ( .I(n1927), .ZN(n1928) );
  and2 U2937 ( .A1(n1931), .A2(n1822), .Z(n1070) );
  and2 U2938 ( .A1(n1835), .A2(n1824), .Z(n1071) );
  and2 U2939 ( .A1(n1833), .A2(n1832), .Z(n1041) );
  and2 U2940 ( .A1(n1835), .A2(n1834), .Z(n1042) );
  and2 U2941 ( .A1(n1010), .A2(n1011), .Z(n997) );
  or2 U2942 ( .A1(n999), .A2(n1000), .Z(n998) );
  or2 U2943 ( .A1(n977), .A2(n978), .Z(n976) );
  or2 U2944 ( .A1(n881), .A2(n882), .Z(n880) );
  and2 U2945 ( .A1(n1749), .A2(n883), .Z(n882) );
  and2 U2946 ( .A1(n842), .A2(n843), .Z(n840) );
  or2 U2947 ( .A1(n1934), .A2(n1933), .Z(n1935) );
  and2 U2948 ( .A1(n1936), .A2(n1952), .Z(n1934) );
  or2 U2949 ( .A1(n1939), .A2(n1938), .Z(n1949) );
  or2 U2950 ( .A1(n650), .A2(n651), .Z(n649) );
  inv1 U2951 ( .I(n1845), .ZN(n651) );
  and2 U2952 ( .A1(n530), .A2(n531), .Z(n522) );
  or2 U2953 ( .A1(n381), .A2(n537), .Z(n530) );
  and2 U2954 ( .A1(n445), .A2(n446), .Z(n443) );
  or2 U2955 ( .A1(n381), .A2(n451), .Z(n445) );
  and2 U2956 ( .A1(n372), .A2(n373), .Z(n370) );
  or2 U2957 ( .A1(n381), .A2(n382), .Z(n372) );
  or2 U2958 ( .A1(n795), .A2(n796), .Z(s5) );
  or2 U2959 ( .A1(n716), .A2(n717), .Z(t5) );
  or2 U2960 ( .A1(n628), .A2(n629), .Z(u5) );
  or2 U2961 ( .A1(n575), .A2(n576), .Z(v5) );
  or2 U2962 ( .A1(n423), .A2(n424), .Z(x5) );
  or2 U2963 ( .A1(n350), .A2(n351), .Z(y5) );
  or2 U2964 ( .A1(n288), .A2(n289), .Z(z5) );
  or2 U2965 ( .A1(n1668), .A2(n1669), .Z(a6) );
  and2 U2966 ( .A1(n1951), .A2(n1852), .Z(c6) );
  and2 U2967 ( .A1(n1857), .A2(n1856), .Z(d6) );
  and2 U2968 ( .A1(n1358), .A2(n1951), .Z(e6) );
  and2 U2969 ( .A1(n1861), .A2(n1862), .Z(f6) );
  and2 U2970 ( .A1(n1865), .A2(n1864), .Z(g6) );
  and2 U2971 ( .A1(n1869), .A2(n1868), .Z(h6) );
  or2 U2972 ( .A1(n948), .A2(n949), .Z(o6) );
  or2 U2973 ( .A1(n910), .A2(n911), .Z(p6) );
  or2 U2974 ( .A1(n874), .A2(n875), .Z(q6) );
  or2 U2975 ( .A1(n1885), .A2(n623), .Z(s6) );
  or2 U2976 ( .A1(n621), .A2(n622), .Z(u6) );
  or2 U2977 ( .A1(n481), .A2(n415), .Z(w6) );
  and2 U2978 ( .A1(n414), .A2(n338), .Z(x6) );
  and2 U2979 ( .A1(n337), .A2(n338), .Z(y6) );
  or2 U2980 ( .A1(n278), .A2(n279), .Z(z6) );
  or2 U2981 ( .A1(n1496), .A2(n1497), .Z(b7) );
  or2 U2982 ( .A1(n1286), .A2(n1287), .Z(f7) );
  or2 U2983 ( .A1(b), .A2(n1113), .Z(i7) );
  or2 U2984 ( .A1(b), .A2(n1109), .Z(j7) );
  or2 U2985 ( .A1(n1060), .A2(b), .Z(k7) );
  or2 U2986 ( .A1(n1031), .A2(n1032), .Z(l7) );
  or2 U2987 ( .A1(n991), .A2(b), .Z(m7) );
  or2 U2988 ( .A1(b), .A2(n971), .Z(n7) );
  or2 U2989 ( .A1(n938), .A2(b), .Z(o7) );
  or2 U2990 ( .A1(n902), .A2(n903), .Z(p7) );
  or2 U2991 ( .A1(n864), .A2(b), .Z(q7) );
  or2 U2992 ( .A1(n831), .A2(n832), .Z(r7) );
  and2 U2993 ( .A1(n613), .A2(n614), .Z(u7) );
  or2 U2994 ( .A1(n475), .A2(n476), .Z(w7) );
  or2 U2995 ( .A1(n1490), .A2(n1491), .Z(b8) );
  and2 U2996 ( .A1(n1427), .A2(n1428), .Z(c8) );
  or2 U2997 ( .A1(n857), .A2(n858), .Z(q8) );
  and2 U2998 ( .A1(n828), .A2(n829), .Z(r8) );
  or2 U2999 ( .A1(n1464), .A2(n1465), .Z(b9) );
  or2 U3000 ( .A1(n1365), .A2(n1366), .Z(d9) );
  or2 U3001 ( .A1(n1156), .A2(n1157), .Z(h9) );
  or2 U3002 ( .A1(n983), .A2(z), .Z(m9) );
  or2 U3003 ( .A1(n954), .A2(n955), .Z(n9) );
  or2 U3004 ( .A1(n919), .A2(z), .Z(o9) );
  or2 U3005 ( .A1(z), .A2(n885), .Z(p9) );
  or2 U3006 ( .A1(n847), .A2(z), .Z(q9) );
  or2 U3007 ( .A1(n820), .A2(n821), .Z(r9) );
  or2 U3008 ( .A1(n761), .A2(z), .Z(s9) );
  or2 U3009 ( .A1(n656), .A2(n657), .Z(t9) );
  and2 U3010 ( .A1(n452), .A2(n453), .Z(w9) );
  and2 U3011 ( .A1(n1954), .A2(n1904), .Z(y9) );
  and2 U3012 ( .A1(n1909), .A2(n1908), .Z(z9) );
  and2 U3013 ( .A1(n1688), .A2(n1954), .Z(a10) );
  and2 U3014 ( .A1(n1913), .A2(n1914), .Z(b10) );
  and2 U3015 ( .A1(n1917), .A2(n1916), .Z(c10) );
  and2 U3016 ( .A1(n1921), .A2(n1920), .Z(d10) );
  or2 U3017 ( .A1(n1070), .A2(n1071), .Z(k10) );
  or2 U3018 ( .A1(n1041), .A2(n1042), .Z(l10) );
  and2 U3019 ( .A1(n997), .A2(n998), .Z(m10) );
  and2 U3020 ( .A1(n976), .A2(n1756), .Z(n10) );
  and2 U3021 ( .A1(n841), .A2(n880), .Z(q10) );
  and2 U3022 ( .A1(n840), .A2(n841), .Z(r10) );
  or2 U3023 ( .A1(n1935), .A2(n650), .Z(s10) );
  or2 U3024 ( .A1(n648), .A2(n649), .Z(u10) );
  or2 U3025 ( .A1(n522), .A2(n444), .Z(w10) );
  and2 U3026 ( .A1(n443), .A2(n371), .Z(x10) );
  and2 U3027 ( .A1(n370), .A2(n371), .Z(y10) );
endmodule

