
module f51m ( x8, x7, x6, x5, x4, x3, x2, x1, x51, x50, x49, x48, x47, x46, 
        x45, x44 );
  input x8, x7, x6, x5, x4, x3, x2, x1;
  output x51, x50, x49, x48, x47, x46, x45, x44;
  wire   n145, n146, n147, n141, n20, n21, n22, n23, n24, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n56, n57, n58, n59,
         n60, n63, n64, n65, n67, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n109, n110, n111, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n129, n130, n131, n132, n133,
         n134, n136, n137, n138, n139, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172;

  or2f U3 ( .A1(n22), .A2(n141), .Z(n21) );
  and2f U4 ( .A1(n23), .A2(n24), .Z(n22) );
  or2f U6 ( .A1(n27), .A2(n28), .Z(n26) );
  or2f U7 ( .A1(n29), .A2(x6), .Z(n23) );
  or2f U9 ( .A1(n147), .A2(n30), .Z(n20) );
  and2f U10 ( .A1(n31), .A2(n32), .Z(n30) );
  or2f U12 ( .A1(n145), .A2(n34), .Z(n33) );
  and2f U13 ( .A1(n35), .A2(n36), .Z(n34) );
  and2f U14 ( .A1(n37), .A2(n38), .Z(n31) );
  and2f U17 ( .A1(x7), .A2(x5), .Z(n39) );
  or2f U30 ( .A1(n57), .A2(n170), .Z(x46) );
  and2f U32 ( .A1(n58), .A2(n148), .Z(n57) );
  or2f U33 ( .A1(n60), .A2(n59), .Z(n58) );
  and2f U36 ( .A1(n145), .A2(n147), .Z(n63) );
  inv1f U38 ( .I(n65), .ZN(n64) );
  and2f U41 ( .A1(n141), .A2(n150), .Z(n65) );
  and2f U47 ( .A1(x3), .A2(n72), .Z(n71) );
  or2f U48 ( .A1(n74), .A2(n73), .Z(n72) );
  or2f U49 ( .A1(n75), .A2(n76), .Z(n74) );
  and2f U50 ( .A1(n51), .A2(n147), .Z(n73) );
  and2f U53 ( .A1(n77), .A2(x5), .Z(n70) );
  or2f U54 ( .A1(n78), .A2(n79), .Z(x45) );
  and2f U65 ( .A1(x5), .A2(x8), .Z(n27) );
  or2f U67 ( .A1(n36), .A2(n95), .Z(n37) );
  or2f U68 ( .A1(n28), .A2(n35), .Z(n95) );
  and2f U71 ( .A1(n96), .A2(x2), .Z(n78) );
  or2f U72 ( .A1(n97), .A2(n98), .Z(n96) );
  or2f U73 ( .A1(n99), .A2(n100), .Z(n98) );
  and2f U75 ( .A1(n102), .A2(n103), .Z(n99) );
  and2f U78 ( .A1(n148), .A2(n147), .Z(n102) );
  or2f U79 ( .A1(n105), .A2(n104), .Z(n97) );
  or2f U80 ( .A1(n77), .A2(n75), .Z(n105) );
  and2f U81 ( .A1(n147), .A2(n169), .Z(n77) );
  or2f U85 ( .A1(n110), .A2(n111), .Z(x44) );
  and2f U88 ( .A1(x1), .A2(n115), .Z(n114) );
  or2f U89 ( .A1(n116), .A2(n117), .Z(n115) );
  or2f U92 ( .A1(n121), .A2(n84), .Z(n119) );
  and2f U96 ( .A1(n123), .A2(n147), .Z(n121) );
  and2f U101 ( .A1(x8), .A2(x7), .Z(n40) );
  or2f U109 ( .A1(n131), .A2(n130), .Z(n129) );
  or2f U110 ( .A1(n75), .A2(n132), .Z(n131) );
  and2f U112 ( .A1(n141), .A2(n134), .Z(n75) );
  buf0 U131 ( .I(n147), .Z(x47) );
  buf0 U132 ( .I(n146), .Z(x50) );
  buf0 U133 ( .I(n145), .Z(x51) );
  and2f U134 ( .A1(n21), .A2(x4), .Z(n168) );
  or2 U135 ( .A1(n80), .A2(n81), .Z(n79) );
  and2 U136 ( .A1(n64), .A2(n160), .Z(n158) );
  or2 U137 ( .A1(n153), .A2(n154), .Z(n111) );
  or2f U138 ( .A1(n27), .A2(n94), .Z(n93) );
  inv1 U139 ( .I(x5), .ZN(n148) );
  and2f U140 ( .A1(n109), .A2(n149), .Z(n104) );
  and2f U141 ( .A1(n141), .A2(x3), .Z(n149) );
  inv1 U142 ( .I(x5), .ZN(n35) );
  or2 U143 ( .A1(n28), .A2(n33), .Z(n32) );
  and2 U144 ( .A1(n133), .A2(n147), .Z(n137) );
  and2 U145 ( .A1(n88), .A2(n89), .Z(n80) );
  and2 U146 ( .A1(n87), .A2(n147), .Z(n88) );
  inv1 U147 ( .I(x8), .ZN(n145) );
  inv1 U148 ( .I(x6), .ZN(n28) );
  or2 U149 ( .A1(n71), .A2(n157), .Z(n170) );
  buf0 U150 ( .I(n40), .Z(n150) );
  inv1 U151 ( .I(x7), .ZN(n36) );
  or2f U152 ( .A1(n137), .A2(n136), .Z(n151) );
  and2 U153 ( .A1(n151), .A2(n152), .Z(n162) );
  and2 U154 ( .A1(n67), .A2(x1), .Z(n152) );
  and2 U155 ( .A1(n119), .A2(n155), .Z(n153) );
  and2f U156 ( .A1(x3), .A2(n114), .Z(n154) );
  and2 U157 ( .A1(n120), .A2(x3), .Z(n155) );
  and2f U158 ( .A1(n69), .A2(n166), .Z(n164) );
  inv1f U159 ( .I(n167), .ZN(n29) );
  and2f U160 ( .A1(n118), .A2(n141), .Z(n116) );
  or2f U161 ( .A1(n64), .A2(x3), .Z(n156) );
  inv1f U162 ( .I(n156), .ZN(n165) );
  or2f U163 ( .A1(n70), .A2(n56), .Z(n157) );
  or2f U164 ( .A1(n159), .A2(n158), .Z(n60) );
  and2f U165 ( .A1(x3), .A2(n63), .Z(n159) );
  and2 U166 ( .A1(n28), .A2(x3), .Z(n160) );
  and2 U167 ( .A1(n129), .A2(n163), .Z(n161) );
  or2f U168 ( .A1(n162), .A2(n161), .Z(n110) );
  and2 U169 ( .A1(n120), .A2(n67), .Z(n163) );
  or2f U170 ( .A1(n165), .A2(n164), .Z(n59) );
  and2 U171 ( .A1(x6), .A2(n67), .Z(n166) );
  or2f U172 ( .A1(n39), .A2(n40), .Z(n167) );
  or2f U173 ( .A1(n167), .A2(n26), .Z(n24) );
  and2f U174 ( .A1(n20), .A2(n168), .Z(n141) );
  and2 U175 ( .A1(n106), .A2(n67), .Z(n169) );
  inv1f U176 ( .I(n141), .ZN(n147) );
  and2 U177 ( .A1(x7), .A2(x8), .Z(n171) );
  or2f U178 ( .A1(n171), .A2(n172), .Z(n38) );
  or2f U179 ( .A1(x6), .A2(n39), .Z(n172) );
  and2 U180 ( .A1(x2), .A2(n141), .Z(n130) );
  or2 U181 ( .A1(n141), .A2(n150), .Z(n69) );
  and2 U182 ( .A1(x3), .A2(n150), .Z(n94) );
  and2 U183 ( .A1(x2), .A2(n124), .Z(n117) );
  and2 U184 ( .A1(n109), .A2(n125), .Z(n124) );
  or2 U185 ( .A1(n150), .A2(x5), .Z(n125) );
  or2 U186 ( .A1(n109), .A2(n122), .Z(n118) );
  or2 U187 ( .A1(x2), .A2(n150), .Z(n122) );
  inv1 U188 ( .I(n133), .ZN(n132) );
  inv1 U189 ( .I(x1), .ZN(n120) );
  or2 U190 ( .A1(n43), .A2(n148), .Z(n86) );
  inv1 U191 ( .I(n118), .ZN(n84) );
  or2 U192 ( .A1(n83), .A2(n84), .Z(n82) );
  and2 U193 ( .A1(n85), .A2(n86), .Z(n83) );
  and2 U194 ( .A1(n87), .A2(n67), .Z(n85) );
  and2 U195 ( .A1(n94), .A2(n101), .Z(n100) );
  or2 U196 ( .A1(n90), .A2(n91), .Z(n89) );
  and2 U197 ( .A1(x3), .A2(x5), .Z(n90) );
  and2 U198 ( .A1(n49), .A2(n148), .Z(n48) );
  or2 U199 ( .A1(n50), .A2(n51), .Z(n49) );
  and2 U200 ( .A1(x5), .A2(n43), .Z(n47) );
  inv1 U201 ( .I(n146), .ZN(n52) );
  and2 U202 ( .A1(n28), .A2(n36), .Z(n43) );
  or2 U203 ( .A1(x7), .A2(n145), .Z(n44) );
  or2 U204 ( .A1(n53), .A2(n50), .Z(n146) );
  or2 U205 ( .A1(n106), .A2(n138), .Z(n133) );
  or2 U206 ( .A1(n148), .A2(n87), .Z(n138) );
  inv1 U207 ( .I(n101), .ZN(n109) );
  and2 U208 ( .A1(n86), .A2(n87), .Z(n136) );
  and2 U209 ( .A1(n148), .A2(n28), .Z(n101) );
  inv1 U210 ( .I(n94), .ZN(n103) );
  inv1 U211 ( .I(x2), .ZN(n87) );
  or2 U212 ( .A1(n76), .A2(n92), .Z(n91) );
  and2 U213 ( .A1(n93), .A2(x6), .Z(n92) );
  or2 U214 ( .A1(n28), .A2(n139), .Z(n106) );
  and2 U215 ( .A1(n36), .A2(n145), .Z(n139) );
  inv1 U216 ( .I(n86), .ZN(n134) );
  inv1 U217 ( .I(n37), .ZN(n76) );
  and2 U218 ( .A1(x6), .A2(n53), .Z(n51) );
  and2 U219 ( .A1(n36), .A2(x8), .Z(n53) );
  and2 U220 ( .A1(x7), .A2(n145), .Z(n50) );
  inv1 U221 ( .I(n117), .ZN(n123) );
  inv1 U222 ( .I(x3), .ZN(n67) );
  and2 U223 ( .A1(n47), .A2(n67), .Z(n56) );
  and2 U224 ( .A1(n82), .A2(n141), .Z(n81) );
  and2 U225 ( .A1(x5), .A2(n52), .Z(n45) );
  or2 U226 ( .A1(n47), .A2(n48), .Z(n46) );
  and2 U227 ( .A1(n44), .A2(x6), .Z(n41) );
  and2 U228 ( .A1(n43), .A2(x8), .Z(n42) );
  or2 U229 ( .A1(n45), .A2(n46), .Z(x48) );
  or2 U230 ( .A1(n41), .A2(n42), .Z(x49) );
endmodule

