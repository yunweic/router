
module example2 ( h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, 
        s1, r1, q1, p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, 
        a1, z0, y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, 
        i0, h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, 
        n, m, l, k, j, i, h, g, f, e, d, b, a, v4, u4, t4, s4, r4, q4, p4, o4, 
        n4, m4, l4, k4, j4, i4, h4, g4, f4, e4, d4, c4, b4, a4, z3, y3, x3, w3, 
        v3, u3, t3, s3, r3, q3, p3, o3, n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, 
        d3, c3, b3, a3, z2, y2, x2, w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, 
        l2, k2, j2, i2 );
  input h2, g2, f2, e2, d2, c2, b2, a2, z1, y1, x1, w1, v1, u1, t1, s1, r1, q1,
         p1, o1, n1, m1, l1, k1, j1, i1, h1, g1, f1, e1, d1, c1, b1, a1, z0,
         y0, x0, w0, v0, u0, t0, s0, r0, q0, p0, o0, n0, m0, l0, k0, j0, i0,
         h0, g0, f0, e0, d0, c0, b0, a0, z, y, x, w, v, u, t, s, r, q, p, o, n,
         m, l, k, j, i, h, g, f, e, d, b, a;
  output v4, u4, t4, s4, r4, q4, p4, o4, n4, m4, l4, k4, j4, i4, h4, g4, f4,
         e4, d4, c4, b4, a4, z3, y3, x3, w3, v3, u3, t3, s3, r3, q3, p3, o3,
         n3, m3, l3, k3, j3, i3, h3, g3, f3, e3, d3, c3, b3, a3, z2, y2, x2,
         w2, v2, u2, t2, s2, r2, q2, p2, o2, n2, m2, l2, k2, j2, i2;
  wire   n323, n324, n325, n6, n7, n9, n10, n11, n12, n13, n14, n16, n17, n18,
         n19, n20, n21, n24, n25, n26, n27, n30, n31, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n65, n69, n71, n72, n73, n74,
         n75, n76, n78, n79, n80, n81, n82, n83, n85, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n108, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n206, n207, n208, n213, n226, n228, n245, n246,
         n247, n248, n249, n250, n251, n252, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n326, n327;

  or2 U2 ( .A1(n6), .A2(n7), .Z(z2) );
  and2 U3 ( .A1(x0), .A2(p0), .Z(n7) );
  and2 U4 ( .A1(k0), .A2(n255), .Z(n6) );
  or2 U6 ( .A1(n9), .A2(n10), .Z(y2) );
  and2 U7 ( .A1(y0), .A2(p0), .Z(n10) );
  and2 U8 ( .A1(j0), .A2(n255), .Z(n9) );
  or2 U10 ( .A1(n11), .A2(n12), .Z(x2) );
  and2 U11 ( .A1(z0), .A2(p0), .Z(n12) );
  and2 U12 ( .A1(i0), .A2(n255), .Z(n11) );
  or2 U14 ( .A1(n13), .A2(n14), .Z(w2) );
  and2 U15 ( .A1(h0), .A2(n255), .Z(n14) );
  and2 U16 ( .A1(a1), .A2(p0), .Z(n13) );
  and2 U17 ( .A1(n315), .A2(h2), .Z(v4) );
  or2 U19 ( .A1(n16), .A2(n17), .Z(v2) );
  and2 U20 ( .A1(g1), .A2(p0), .Z(n17) );
  and2 U21 ( .A1(g0), .A2(n255), .Z(n16) );
  or2 U22 ( .A1(n18), .A2(n19), .Z(u4) );
  and2 U24 ( .A1(n20), .A2(n21), .Z(n18) );
  and2 U25 ( .A1(n320), .A2(n322), .Z(n21) );
  or2 U27 ( .A1(n24), .A2(n25), .Z(u2) );
  and2 U28 ( .A1(h1), .A2(p0), .Z(n25) );
  and2 U29 ( .A1(f0), .A2(n255), .Z(n24) );
  and2 U30 ( .A1(n315), .A2(f2), .Z(t4) );
  or2 U32 ( .A1(n26), .A2(n27), .Z(t2) );
  and2 U33 ( .A1(i1), .A2(p0), .Z(n27) );
  and2 U34 ( .A1(e0), .A2(n255), .Z(n26) );
  or2 U38 ( .A1(n30), .A2(n31), .Z(s2) );
  and2 U39 ( .A1(j1), .A2(p0), .Z(n31) );
  and2 U40 ( .A1(d0), .A2(n255), .Z(n30) );
  and2 U41 ( .A1(n315), .A2(d2), .Z(r4) );
  and2 U44 ( .A1(n36), .A2(n317), .Z(n35) );
  or2 U47 ( .A1(n40), .A2(n41), .Z(r2) );
  and2 U48 ( .A1(p0), .A2(k1), .Z(n41) );
  and2 U49 ( .A1(c0), .A2(n255), .Z(n40) );
  or2 U50 ( .A1(n42), .A2(n43), .Z(q4) );
  and2 U51 ( .A1(n44), .A2(n322), .Z(n43) );
  or2 U52 ( .A1(n45), .A2(n46), .Z(n44) );
  or2 U53 ( .A1(n47), .A2(n48), .Z(n46) );
  and2 U54 ( .A1(n39), .A2(n49), .Z(n48) );
  and2 U55 ( .A1(n50), .A2(n49), .Z(n42) );
  or2 U57 ( .A1(n51), .A2(n52), .Z(q2) );
  and2 U58 ( .A1(l1), .A2(p0), .Z(n52) );
  and2 U59 ( .A1(b0), .A2(n255), .Z(n51) );
  and2 U60 ( .A1(n53), .A2(n322), .Z(p4) );
  or2 U61 ( .A1(n45), .A2(n54), .Z(n53) );
  or2 U62 ( .A1(n55), .A2(n56), .Z(n54) );
  and2 U63 ( .A1(n47), .A2(a2), .Z(n56) );
  and2 U64 ( .A1(p0), .A2(n57), .Z(n55) );
  or2 U65 ( .A1(n58), .A2(n59), .Z(n57) );
  and2 U66 ( .A1(a2), .A2(n60), .Z(n58) );
  or2 U67 ( .A1(n61), .A2(n62), .Z(n45) );
  and2 U73 ( .A1(g), .A2(r0), .Z(n69) );
  or2 U74 ( .A1(n71), .A2(n72), .Z(p2) );
  and2 U75 ( .A1(m1), .A2(p0), .Z(n72) );
  and2 U76 ( .A1(a0), .A2(n255), .Z(n71) );
  and2 U78 ( .A1(n75), .A2(n76), .Z(n74) );
  or2 U79 ( .A1(n321), .A2(n78), .Z(n76) );
  or2 U80 ( .A1(n39), .A2(n79), .Z(n78) );
  and2 U81 ( .A1(n80), .A2(n38), .Z(n79) );
  and2 U82 ( .A1(p0), .A2(n65), .Z(n80) );
  and2 U83 ( .A1(n322), .A2(n60), .Z(n75) );
  and2 U84 ( .A1(n81), .A2(n59), .Z(n73) );
  and2 U86 ( .A1(n318), .A2(n83), .Z(n81) );
  and2 U88 ( .A1(r0), .A2(n255), .Z(n85) );
  inv1 U90 ( .I(r0), .ZN(n65) );
  or2 U92 ( .A1(n87), .A2(n88), .Z(o2) );
  and2 U93 ( .A1(z), .A2(n255), .Z(n88) );
  and2 U94 ( .A1(n1), .A2(p0), .Z(n87) );
  and2 U95 ( .A1(n89), .A2(n90), .Z(n4) );
  inv1 U96 ( .I(n91), .ZN(n90) );
  or2 U97 ( .A1(b), .A2(d), .Z(n91) );
  and2 U98 ( .A1(e), .A2(a), .Z(n89) );
  or2 U100 ( .A1(n92), .A2(n93), .Z(n2) );
  and2 U101 ( .A1(y), .A2(n255), .Z(n93) );
  and2 U102 ( .A1(o1), .A2(p0), .Z(n92) );
  or2 U103 ( .A1(n94), .A2(n95), .Z(m4) );
  or2 U104 ( .A1(n96), .A2(n97), .Z(n95) );
  or2 U105 ( .A1(b), .A2(n98), .Z(n94) );
  and2 U106 ( .A1(n99), .A2(c2), .Z(n98) );
  and2 U107 ( .A1(n100), .A2(n101), .Z(n99) );
  or2 U108 ( .A1(z1), .A2(n49), .Z(n100) );
  and2 U114 ( .A1(g2), .A2(h2), .Z(n108) );
  or2 U116 ( .A1(n110), .A2(n111), .Z(k4) );
  and2 U117 ( .A1(p), .A2(n112), .Z(n111) );
  and2 U118 ( .A1(x), .A2(n326), .Z(n110) );
  or2 U120 ( .A1(n114), .A2(n115), .Z(j4) );
  or2 U121 ( .A1(n116), .A2(n117), .Z(n115) );
  and2 U122 ( .A1(w), .A2(n326), .Z(n117) );
  and2 U123 ( .A1(w1), .A2(n118), .Z(n116) );
  and2 U124 ( .A1(o), .A2(n112), .Z(n114) );
  and2 U126 ( .A1(n119), .A2(n322), .Z(j2) );
  or2 U127 ( .A1(n60), .A2(n120), .Z(n119) );
  or2 U128 ( .A1(n82), .A2(n96), .Z(n120) );
  and2 U129 ( .A1(n320), .A2(n319), .Z(n96) );
  or2 U130 ( .A1(n122), .A2(n123), .Z(i4) );
  or2 U131 ( .A1(n124), .A2(n125), .Z(n123) );
  and2 U132 ( .A1(v), .A2(n327), .Z(n125) );
  and2 U133 ( .A1(v1), .A2(n118), .Z(n124) );
  and2 U134 ( .A1(n), .A2(n112), .Z(n122) );
  or2 U136 ( .A1(n126), .A2(n127), .Z(i2) );
  and2 U137 ( .A1(h), .A2(n255), .Z(n127) );
  and2 U138 ( .A1(p0), .A2(n128), .Z(n126) );
  or2 U139 ( .A1(b1), .A2(n323), .Z(n128) );
  or2 U140 ( .A1(n129), .A2(n318), .Z(n323) );
  and2 U141 ( .A1(n101), .A2(n322), .Z(n129) );
  inv1 U142 ( .I(n82), .ZN(n101) );
  or2 U143 ( .A1(n130), .A2(n131), .Z(h4) );
  or2 U144 ( .A1(n132), .A2(n133), .Z(n131) );
  and2 U145 ( .A1(u), .A2(n113), .Z(n133) );
  and2 U146 ( .A1(u1), .A2(n118), .Z(n132) );
  and2 U147 ( .A1(m), .A2(n112), .Z(n130) );
  or2 U149 ( .A1(n134), .A2(n135), .Z(g4) );
  or2 U150 ( .A1(n136), .A2(n137), .Z(n135) );
  and2 U151 ( .A1(t), .A2(n113), .Z(n137) );
  and2 U152 ( .A1(t1), .A2(n118), .Z(n136) );
  and2 U153 ( .A1(l), .A2(n112), .Z(n134) );
  and2 U154 ( .A1(n138), .A2(n139), .Z(g3) );
  and2 U155 ( .A1(n322), .A2(n140), .Z(n139) );
  and2 U156 ( .A1(g), .A2(n141), .Z(n138) );
  or2 U157 ( .A1(n62), .A2(n316), .Z(n141) );
  or2 U158 ( .A1(n142), .A2(n143), .Z(f4) );
  or2 U159 ( .A1(n144), .A2(n145), .Z(n143) );
  and2 U160 ( .A1(s), .A2(n326), .Z(n145) );
  and2 U161 ( .A1(s1), .A2(n118), .Z(n144) );
  and2 U162 ( .A1(k), .A2(n112), .Z(n142) );
  or2 U163 ( .A1(n97), .A2(n146), .Z(f3) );
  or2 U164 ( .A1(b), .A2(n147), .Z(n146) );
  and2 U165 ( .A1(n62), .A2(g), .Z(n147) );
  and2 U166 ( .A1(n321), .A2(n60), .Z(n62) );
  inv1 U167 ( .I(a), .ZN(n97) );
  or2 U168 ( .A1(n148), .A2(n149), .Z(e4) );
  or2 U169 ( .A1(n150), .A2(n151), .Z(n149) );
  and2 U170 ( .A1(r), .A2(n327), .Z(n151) );
  and2 U171 ( .A1(r1), .A2(n118), .Z(n150) );
  and2 U172 ( .A1(j), .A2(n112), .Z(n148) );
  and2 U194 ( .A1(p1), .A2(n50), .Z(n168) );
  and2 U195 ( .A1(n169), .A2(y1), .Z(n167) );
  and2 U196 ( .A1(n39), .A2(n318), .Z(n169) );
  or2 U198 ( .A1(n170), .A2(n171), .Z(d4) );
  or2 U199 ( .A1(n172), .A2(n173), .Z(n171) );
  and2 U200 ( .A1(q), .A2(n113), .Z(n173) );
  and2 U202 ( .A1(n320), .A2(f), .Z(n174) );
  and2 U204 ( .A1(n322), .A2(n47), .Z(n175) );
  and2 U205 ( .A1(n118), .A2(n176), .Z(n172) );
  or2 U206 ( .A1(q1), .A2(y1), .Z(n176) );
  and2 U207 ( .A1(n317), .A2(n50), .Z(n118) );
  and2 U209 ( .A1(n319), .A2(a2), .Z(n38) );
  and2 U215 ( .A1(i), .A2(n112), .Z(n170) );
  and2 U216 ( .A1(n179), .A2(n20), .Z(n112) );
  and2 U217 ( .A1(n47), .A2(f), .Z(n20) );
  inv1 U219 ( .I(c2), .ZN(n60) );
  and2 U220 ( .A1(n320), .A2(n180), .Z(n179) );
  and2 U221 ( .A1(n181), .A2(n322), .Z(n180) );
  inv1 U222 ( .I(b1), .ZN(n181) );
  or2 U224 ( .A1(n182), .A2(n183), .Z(d3) );
  and2 U225 ( .A1(t0), .A2(p0), .Z(n183) );
  and2 U226 ( .A1(o0), .A2(n255), .Z(n182) );
  or2 U228 ( .A1(n184), .A2(n185), .Z(c3) );
  and2 U229 ( .A1(u0), .A2(p0), .Z(n185) );
  and2 U230 ( .A1(n0), .A2(n255), .Z(n184) );
  or2 U232 ( .A1(n186), .A2(n187), .Z(b3) );
  and2 U233 ( .A1(v0), .A2(p0), .Z(n187) );
  and2 U234 ( .A1(m0), .A2(n255), .Z(n186) );
  or2 U266 ( .A1(n206), .A2(n207), .Z(a3) );
  and2 U267 ( .A1(w0), .A2(p0), .Z(n207) );
  and2 U268 ( .A1(l0), .A2(n255), .Z(n206) );
  and2 U270 ( .A1(n251), .A2(e2), .Z(n208) );
  and2 U272 ( .A1(n213), .A2(g), .Z(h3) );
  and2 U274 ( .A1(n213), .A2(t0), .Z(i3) );
  inv1 U275 ( .I(n247), .ZN(n213) );
  and2 U276 ( .A1(n213), .A2(u0), .Z(j3) );
  and2 U278 ( .A1(n213), .A2(v0), .Z(k3) );
  and2 U279 ( .A1(n213), .A2(w0), .Z(l3) );
  and2 U280 ( .A1(n213), .A2(x0), .Z(m3) );
  and2 U281 ( .A1(n213), .A2(y0), .Z(n3) );
  and2 U282 ( .A1(n213), .A2(z0), .Z(o3) );
  buf0 U304 ( .I(n325), .Z(k2) );
  buf0 U305 ( .I(n324), .Z(l2) );
  buf0 U306 ( .I(n323), .Z(m2) );
  or2 U309 ( .A1(n283), .A2(r0), .Z(n247) );
  or2 U312 ( .A1(n247), .A2(n250), .Z(n249) );
  inv1 U313 ( .I(n249), .ZN(n297) );
  inv1 U314 ( .I(a1), .ZN(n250) );
  inv1 U315 ( .I(f2), .ZN(n251) );
  or2 U316 ( .A1(n245), .A2(n208), .Z(n252) );
  inv1 U319 ( .I(p0), .ZN(n255) );
  inv1 U320 ( .I(b), .ZN(n322) );
  inv1 U322 ( .I(b2), .ZN(n319) );
  inv1 U325 ( .I(e2), .ZN(n307) );
  and2 U326 ( .A1(n307), .A2(h2), .Z(n257) );
  inv1 U330 ( .I(n49), .ZN(n317) );
  inv1 U331 ( .I(f), .ZN(n321) );
  or2 U334 ( .A1(n140), .A2(x1), .Z(n258) );
  or2 U335 ( .A1(n258), .A2(g2), .Z(n262) );
  inv1 U336 ( .I(d2), .ZN(n306) );
  or2 U337 ( .A1(n307), .A2(n306), .Z(n260) );
  inv1 U338 ( .I(f2), .ZN(n308) );
  or2 U339 ( .A1(n285), .A2(n308), .Z(n259) );
  and2 U343 ( .A1(n65), .A2(n268), .Z(n263) );
  or2 U344 ( .A1(n263), .A2(n85), .Z(n83) );
  and2 U345 ( .A1(n59), .A2(n65), .Z(n264) );
  and2 U346 ( .A1(n265), .A2(n264), .Z(n61) );
  inv1 U347 ( .I(n35), .ZN(n266) );
  inv1 U348 ( .I(n316), .ZN(n281) );
  and2 U349 ( .A1(n266), .A2(n281), .Z(n267) );
  or2 U352 ( .A1(n168), .A2(n167), .Z(n325) );
  or2 U356 ( .A1(n271), .A2(b), .Z(n273) );
  or2 U357 ( .A1(n319), .A2(n321), .Z(n272) );
  inv1 U359 ( .I(q0), .ZN(n275) );
  and2 U360 ( .A1(n325), .A2(n317), .Z(n274) );
  and2 U361 ( .A1(n275), .A2(n274), .Z(n276) );
  or2 U362 ( .A1(n313), .A2(n276), .Z(e3) );
  inv1 U365 ( .I(n291), .ZN(n288) );
  or2 U366 ( .A1(n288), .A2(h2), .Z(n279) );
  or2 U371 ( .A1(n283), .A2(r0), .Z(n301) );
  inv1 U372 ( .I(g2), .ZN(n284) );
  and2 U373 ( .A1(n284), .A2(h2), .Z(n287) );
  and2 U376 ( .A1(n288), .A2(n289), .Z(n293) );
  inv1 U380 ( .I(n304), .ZN(n294) );
  and2 U381 ( .A1(n294), .A2(n69), .Z(n295) );
  and2 U382 ( .A1(n298), .A2(n295), .Z(n296) );
  or2 U383 ( .A1(n297), .A2(n296), .Z(p3) );
  or2 U384 ( .A1(n304), .A2(n65), .Z(n300) );
  or2 U386 ( .A1(n300), .A2(n299), .Z(n302) );
  and2 U387 ( .A1(n108), .A2(n294), .Z(n305) );
  and2 U388 ( .A1(n306), .A2(n305), .Z(n310) );
  and2 U389 ( .A1(n308), .A2(n307), .Z(n309) );
  and2 U390 ( .A1(n310), .A2(n309), .Z(l4) );
  and2 U391 ( .A1(n315), .A2(e2), .Z(n314) );
  inv1 U392 ( .I(n312), .ZN(n313) );
  or2 U393 ( .A1(n314), .A2(n313), .Z(s4) );
  inv1f U271 ( .I(n248), .ZN(n228) );
  and2f U273 ( .A1(n226), .A2(b1), .Z(q3) );
  and2f U277 ( .A1(n226), .A2(l1), .Z(a4) );
  and2f U283 ( .A1(n226), .A2(f1), .Z(u3) );
  and2f U284 ( .A1(n226), .A2(h1), .Z(w3) );
  and2f U285 ( .A1(n226), .A2(n1), .Z(c4) );
  and2f U286 ( .A1(n226), .A2(k1), .Z(z3) );
  and2f U287 ( .A1(n228), .A2(g1), .Z(v3) );
  and2f U288 ( .A1(n228), .A2(j1), .Z(y3) );
  and2f U289 ( .A1(n228), .A2(m1), .Z(b4) );
  and2f U290 ( .A1(n228), .A2(d1), .Z(s3) );
  and2f U291 ( .A1(n228), .A2(e1), .Z(t3) );
  and2f U292 ( .A1(n228), .A2(i1), .Z(x3) );
  and2f U293 ( .A1(n228), .A2(c1), .Z(r3) );
  or2 U294 ( .A1(n281), .A2(n280), .Z(n304) );
  and2 U295 ( .A1(n82), .A2(n321), .Z(n316) );
  or2 U296 ( .A1(n293), .A2(n292), .Z(n298) );
  or2f U297 ( .A1(n273), .A2(n272), .Z(n312) );
  or2f U298 ( .A1(n73), .A2(n74), .Z(o4) );
  and2 U299 ( .A1(n324), .A2(n174), .Z(n113) );
  and2 U300 ( .A1(n324), .A2(n174), .Z(n327) );
  and2f U301 ( .A1(b1), .A2(n175), .Z(n324) );
  inv1 U302 ( .I(e2), .ZN(n246) );
  inv1 U303 ( .I(a2), .ZN(n320) );
  inv1 U307 ( .I(n265), .ZN(n268) );
  inv1 U308 ( .I(s0), .ZN(n140) );
  inv1 U310 ( .I(n289), .ZN(n290) );
  and2 U311 ( .A1(n324), .A2(n174), .Z(n326) );
  and2 U317 ( .A1(e2), .A2(n285), .Z(n256) );
  and2 U318 ( .A1(n315), .A2(g2), .Z(n19) );
  and2f U321 ( .A1(n318), .A2(n38), .Z(n50) );
  or2 U323 ( .A1(n38), .A2(n39), .Z(n36) );
  inv1f U324 ( .I(n311), .ZN(n315) );
  or2f U327 ( .A1(n257), .A2(n256), .Z(n49) );
  and2f U328 ( .A1(n252), .A2(n290), .Z(n292) );
  or2f U329 ( .A1(n287), .A2(n286), .Z(n289) );
  inv1f U332 ( .I(h2), .ZN(n285) );
  inv1 U333 ( .I(n248), .ZN(n226) );
  and2f U340 ( .A1(a2), .A2(b2), .Z(n82) );
  and2f U341 ( .A1(n82), .A2(f), .Z(n59) );
  or2f U342 ( .A1(n267), .A2(n280), .Z(n311) );
  inv1f U350 ( .I(n280), .ZN(n318) );
  and2f U351 ( .A1(n60), .A2(b2), .Z(n47) );
  or2f U353 ( .A1(b), .A2(n60), .Z(n280) );
  and2f U354 ( .A1(n320), .A2(b2), .Z(n39) );
  or2f U355 ( .A1(n268), .A2(n320), .Z(n269) );
  inv1f U358 ( .I(n298), .ZN(n299) );
  or2f U363 ( .A1(n252), .A2(n285), .Z(n278) );
  and2f U364 ( .A1(g2), .A2(n285), .Z(n286) );
  and2f U367 ( .A1(c2), .A2(n270), .Z(n271) );
  or2f U368 ( .A1(n269), .A2(r0), .Z(n270) );
  or2f U369 ( .A1(n262), .A2(n261), .Z(n265) );
  or2f U370 ( .A1(n260), .A2(n259), .Z(n261) );
  or2f U374 ( .A1(n245), .A2(n277), .Z(n291) );
  and2f U375 ( .A1(n251), .A2(e2), .Z(n277) );
  or2f U377 ( .A1(n282), .A2(n304), .Z(n283) );
  and2f U378 ( .A1(n279), .A2(n278), .Z(n282) );
  and2f U379 ( .A1(f2), .A2(n246), .Z(n245) );
  and2f U385 ( .A1(n301), .A2(n302), .Z(n248) );
endmodule

