
module dalu ( sh0, sh1, sh2, musel1, musel2, musel3, musel4, opsel0, opsel1, 
        opsel2, opsel3, inD0, inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, 
        inD9, inD10, inD11, inD12, inD13, inD14, inD15, inC0, inC1, inC2, inC3, 
        inC4, inC5, inC6, inC7, inC8, inC9, inC10, inC11, inC12, inC13, inC14, 
        inC15, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7, inB8, inB9, 
        inB10, inB11, inB12, inB13, inB14, inB15, inA0, inA1, inA2, inA3, inA4, 
        inA5, inA6, inA7, inA8, inA9, inA10, inA11, inA12, inA13, inA14, inA15, 
        O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15
 );
  input sh0, sh1, sh2, musel1, musel2, musel3, musel4, opsel0, opsel1, opsel2,
         opsel3, inD0, inD1, inD2, inD3, inD4, inD5, inD6, inD7, inD8, inD9,
         inD10, inD11, inD12, inD13, inD14, inD15, inC0, inC1, inC2, inC3,
         inC4, inC5, inC6, inC7, inC8, inC9, inC10, inC11, inC12, inC13, inC14,
         inC15, inB0, inB1, inB2, inB3, inB4, inB5, inB6, inB7, inB8, inB9,
         inB10, inB11, inB12, inB13, inB14, inB15, inA0, inA1, inA2, inA3,
         inA4, inA5, inA6, inA7, inA8, inA9, inA10, inA11, inA12, inA13, inA14,
         inA15;
  output O0, O1, O2, O3, O4, O5, O6, O7, O8, O9, O10, O11, O12, O13, O14, O15;
  wire   n54, n55, n56, n57, n58, n59, n60, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n81, n82, n83,
         n85, n86, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n459, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n487, n488, n489, n490, n491, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952;

  and2f U3 ( .A1(n58), .A2(n59), .Z(n57) );
  and2f U25 ( .A1(n95), .A2(n96), .Z(n94) );
  or2f U26 ( .A1(n97), .A2(n98), .Z(n95) );
  and2f U27 ( .A1(sh0), .A2(n99), .Z(n97) );
  or2f U28 ( .A1(n100), .A2(n101), .Z(n99) );
  and2f U30 ( .A1(n104), .A2(n105), .Z(n93) );
  or2f U31 ( .A1(n106), .A2(n930), .Z(n104) );
  and2f U41 ( .A1(sh2), .A2(n125), .Z(n124) );
  or2f U66 ( .A1(n155), .A2(n156), .Z(n154) );
  and2f U85 ( .A1(n89), .A2(n176), .Z(n155) );
  or2f U86 ( .A1(n177), .A2(n178), .Z(n176) );
  inv1f U87 ( .I(n179), .ZN(n178) );
  and2f U90 ( .A1(n182), .A2(n183), .Z(n181) );
  and2f U93 ( .A1(n186), .A2(n131), .Z(n185) );
  or2f U96 ( .A1(n123), .A2(n190), .Z(n189) );
  and2f U97 ( .A1(sh2), .A2(n102), .Z(n190) );
  or2f U98 ( .A1(n191), .A2(n98), .Z(n186) );
  and2f U99 ( .A1(sh0), .A2(n192), .Z(n191) );
  or2f U100 ( .A1(n193), .A2(n194), .Z(n192) );
  and2f U101 ( .A1(n195), .A2(n196), .Z(n184) );
  or2f U102 ( .A1(n197), .A2(n930), .Z(n195) );
  and2f U106 ( .A1(n58), .A2(n203), .Z(n202) );
  or2f U107 ( .A1(n204), .A2(n205), .Z(n203) );
  and2f U108 ( .A1(n62), .A2(n206), .Z(n205) );
  or2f U131 ( .A1(n229), .A2(n230), .Z(n206) );
  and2f U132 ( .A1(n231), .A2(n196), .Z(n230) );
  or2f U133 ( .A1(n119), .A2(n232), .Z(n196) );
  or2f U134 ( .A1(n233), .A2(n234), .Z(n232) );
  or2f U135 ( .A1(n123), .A2(n235), .Z(n234) );
  or2f U139 ( .A1(n121), .A2(n238), .Z(n237) );
  and2f U140 ( .A1(n198), .A2(n902), .Z(n121) );
  and2f U141 ( .A1(n239), .A2(n240), .Z(n229) );
  and2f U148 ( .A1(n58), .A2(n252), .Z(n251) );
  or2f U149 ( .A1(n253), .A2(n254), .Z(n252) );
  and2f U150 ( .A1(n62), .A2(n255), .Z(n254) );
  or2f U173 ( .A1(n278), .A2(n279), .Z(n255) );
  and2f U174 ( .A1(n280), .A2(n239), .Z(n279) );
  or2f U177 ( .A1(n123), .A2(n284), .Z(n283) );
  or2f U180 ( .A1(n188), .A2(n287), .Z(n286) );
  and2f U181 ( .A1(n247), .A2(n902), .Z(n188) );
  and2f U182 ( .A1(n288), .A2(n289), .Z(n278) );
  or2f U194 ( .A1(n123), .A2(n101), .Z(n304) );
  and2f U195 ( .A1(sh2), .A2(n198), .Z(n101) );
  and2f U226 ( .A1(n58), .A2(n338), .Z(n337) );
  or2f U227 ( .A1(n339), .A2(n340), .Z(n338) );
  and2f U228 ( .A1(n62), .A2(n341), .Z(n340) );
  or2f U251 ( .A1(n365), .A2(n366), .Z(n341) );
  and2f U252 ( .A1(n367), .A2(n308), .Z(n366) );
  or2f U255 ( .A1(n123), .A2(n370), .Z(n369) );
  and2f U256 ( .A1(sh2), .A2(n247), .Z(n129) );
  and2f U260 ( .A1(sh2), .A2(n374), .Z(n373) );
  and2f U261 ( .A1(n313), .A2(n902), .Z(n282) );
  and2f U262 ( .A1(n375), .A2(n376), .Z(n365) );
  and2f U269 ( .A1(n58), .A2(n385), .Z(n384) );
  or2f U270 ( .A1(n386), .A2(n387), .Z(n385) );
  and2f U271 ( .A1(n62), .A2(n388), .Z(n387) );
  or2f U295 ( .A1(n411), .A2(n412), .Z(n388) );
  and2f U296 ( .A1(n413), .A2(n375), .Z(n412) );
  or2f U299 ( .A1(n123), .A2(n193), .Z(n416) );
  and2f U300 ( .A1(sh2), .A2(n293), .Z(n193) );
  or2f U301 ( .A1(n417), .A2(n418), .Z(n293) );
  or2f U306 ( .A1(n422), .A2(n303), .Z(n421) );
  and2f U307 ( .A1(n380), .A2(n902), .Z(n303) );
  and2f U308 ( .A1(sh2), .A2(n423), .Z(n422) );
  and2f U309 ( .A1(n424), .A2(n425), .Z(n411) );
  or2f U314 ( .A1(n430), .A2(n431), .Z(O15) );
  or2f U315 ( .A1(n432), .A2(n433), .Z(n431) );
  and2f U334 ( .A1(n453), .A2(n454), .Z(n432) );
  or2f U360 ( .A1(n936), .A2(n483), .Z(n482) );
  and2f U397 ( .A1(n89), .A2(n525), .Z(n504) );
  or2f U398 ( .A1(n526), .A2(n925), .Z(n525) );
  or2f U422 ( .A1(n551), .A2(n926), .Z(O12) );
  and2f U440 ( .A1(n570), .A2(n136), .Z(n551) );
  or2f U445 ( .A1(n577), .A2(n578), .Z(n570) );
  and2f U447 ( .A1(n952), .A2(n531), .Z(n577) );
  or2f U449 ( .A1(n581), .A2(n582), .Z(n579) );
  or2f U450 ( .A1(n180), .A2(n948), .Z(n582) );
  or2f U459 ( .A1(n226), .A2(n589), .Z(n581) );
  or2f U460 ( .A1(n276), .A2(n227), .Z(n589) );
  and2f U514 ( .A1(n58), .A2(n633), .Z(n632) );
  or2f U535 ( .A1(n654), .A2(n655), .Z(n636) );
  or2f U543 ( .A1(n659), .A2(n660), .Z(n654) );
  and2f U552 ( .A1(n58), .A2(n668), .Z(n667) );
  or2f U553 ( .A1(n669), .A2(n670), .Z(n668) );
  and2f U554 ( .A1(n62), .A2(n671), .Z(n670) );
  or2f U576 ( .A1(n692), .A2(n693), .Z(n277) );
  or2f U577 ( .A1(n361), .A2(n917), .Z(n693) );
  and2f U578 ( .A1(n694), .A2(n695), .Z(n361) );
  and2f U582 ( .A1(n698), .A2(n494), .Z(n697) );
  or2f U586 ( .A1(n408), .A2(n700), .Z(n692) );
  or2f U587 ( .A1(n409), .A2(n701), .Z(n700) );
  and2f U592 ( .A1(n706), .A2(n494), .Z(n705) );
  and2f U605 ( .A1(n688), .A2(n90), .Z(n714) );
  or2f U631 ( .A1(n733), .A2(n734), .Z(n671) );
  and2f U632 ( .A1(n735), .A2(n736), .Z(n734) );
  or2f U642 ( .A1(n284), .A2(n743), .Z(n742) );
  and2f U643 ( .A1(n125), .A2(n902), .Z(n743) );
  or2f U644 ( .A1(n744), .A2(n745), .Z(n125) );
  and2f U647 ( .A1(sh2), .A2(n133), .Z(n284) );
  or2f U649 ( .A1(n119), .A2(n747), .Z(n96) );
  or2f U650 ( .A1(n194), .A2(n748), .Z(n747) );
  or2f U651 ( .A1(n123), .A2(n749), .Z(n748) );
  and2f U652 ( .A1(sh2), .A2(n246), .Z(n749) );
  or2f U653 ( .A1(n750), .A2(n751), .Z(n246) );
  or2f U657 ( .A1(n752), .A2(n753), .Z(n133) );
  or2f U660 ( .A1(n754), .A2(n107), .Z(n746) );
  or2f U662 ( .A1(n547), .A2(n558), .Z(n755) );
  and2f U663 ( .A1(n437), .A2(sh2), .Z(n558) );
  and2f U669 ( .A1(inD12), .A2(n919), .Z(n759) );
  and2f U673 ( .A1(n58), .A2(n764), .Z(n763) );
  or2f U674 ( .A1(n765), .A2(n766), .Z(n764) );
  and2f U675 ( .A1(n62), .A2(n767), .Z(n766) );
  and2f U698 ( .A1(n788), .A2(n789), .Z(n409) );
  and2f U700 ( .A1(n791), .A2(n910), .Z(n790) );
  or2f U701 ( .A1(n917), .A2(n791), .Z(n788) );
  or2f U703 ( .A1(n793), .A2(n782), .Z(n792) );
  or2f U707 ( .A1(n794), .A2(n795), .Z(n767) );
  and2f U708 ( .A1(n796), .A2(n424), .Z(n795) );
  or2f U711 ( .A1(n123), .A2(n238), .Z(n799) );
  and2f U712 ( .A1(sh2), .A2(n313), .Z(n238) );
  or2f U713 ( .A1(n800), .A2(n801), .Z(n313) );
  and2f U714 ( .A1(inD6), .A2(n70), .Z(n801) );
  and2f U720 ( .A1(sh2), .A2(n805), .Z(n804) );
  and2f U721 ( .A1(n429), .A2(n902), .Z(n370) );
  and2f U722 ( .A1(n806), .A2(n807), .Z(n794) );
  or2f U726 ( .A1(n811), .A2(n812), .Z(n198) );
  or2f U770 ( .A1(n852), .A2(n853), .Z(n429) );
  and2f U771 ( .A1(inD4), .A2(n70), .Z(n853) );
  or2f U777 ( .A1(n857), .A2(n858), .Z(n247) );
  and2f U792 ( .A1(n805), .A2(n902), .Z(n864) );
  or2f U793 ( .A1(n865), .A2(n866), .Z(n805) );
  and2f U797 ( .A1(sh2), .A2(n380), .Z(n287) );
  or2f U798 ( .A1(n867), .A2(n868), .Z(n380) );
  or2f U809 ( .A1(n872), .A2(n873), .Z(n374) );
  and2f U816 ( .A1(n828), .A2(n72), .Z(n877) );
  and2f U818 ( .A1(n878), .A2(n494), .Z(n876) );
  and2f U822 ( .A1(n832), .A2(musel3), .Z(n72) );
  and2f U836 ( .A1(n889), .A2(n888), .Z(n701) );
  and2f U838 ( .A1(n891), .A2(n909), .Z(n890) );
  or2f U839 ( .A1(n916), .A2(n891), .Z(n888) );
  or2f U841 ( .A1(n893), .A2(n838), .Z(n892) );
  and2f U846 ( .A1(n900), .A2(musel4), .Z(n494) );
  or2f U848 ( .A1(n452), .A2(n895), .Z(n894) );
  and2f U850 ( .A1(n931), .A2(musel1), .Z(n496) );
  and2f U852 ( .A1(n912), .A2(inC15), .Z(n895) );
  and2f U853 ( .A1(n879), .A2(musel2), .Z(n497) );
  inv1f U854 ( .I(musel1), .ZN(n879) );
  or2f U863 ( .A1(n876), .A2(n877), .Z(n70) );
  and2f U864 ( .A1(n881), .A2(n72), .Z(n419) );
  or2f U865 ( .A1(n876), .A2(n877), .Z(n918) );
  and2 U866 ( .A1(inD13), .A2(n918), .Z(n745) );
  or2 U867 ( .A1(n707), .A2(n394), .Z(n706) );
  and2 U868 ( .A1(inD3), .A2(n919), .Z(n873) );
  and2 U869 ( .A1(inD14), .A2(n919), .Z(n751) );
  or2 U870 ( .A1(n123), .A2(n124), .Z(n122) );
  or2 U871 ( .A1(n119), .A2(n187), .Z(n131) );
  or2 U872 ( .A1(n188), .A2(n189), .Z(n187) );
  or2 U873 ( .A1(n656), .A2(n657), .Z(n655) );
  and2 U874 ( .A1(n496), .A2(inA15), .Z(n452) );
  and2 U875 ( .A1(inD7), .A2(n70), .Z(n418) );
  inv1 U876 ( .I(musel4), .ZN(n832) );
  and2 U877 ( .A1(n293), .A2(n902), .Z(n235) );
  and2 U878 ( .A1(inD5), .A2(n70), .Z(n868) );
  or2 U879 ( .A1(n699), .A2(n347), .Z(n698) );
  and2 U880 ( .A1(inD10), .A2(n70), .Z(n753) );
  inv1 U881 ( .I(n890), .ZN(n889) );
  and2 U882 ( .A1(inD1), .A2(n70), .Z(n866) );
  and2 U883 ( .A1(n374), .A2(n902), .Z(n415) );
  or2 U884 ( .A1(n859), .A2(n860), .Z(n423) );
  and2 U885 ( .A1(inD2), .A2(n919), .Z(n860) );
  and2 U886 ( .A1(inD8), .A2(n70), .Z(n858) );
  or2 U887 ( .A1(n874), .A2(n875), .Z(n851) );
  and2 U888 ( .A1(inD0), .A2(n70), .Z(n875) );
  and2 U889 ( .A1(sh2), .A2(n429), .Z(n307) );
  and2 U890 ( .A1(n944), .A2(n530), .Z(n945) );
  and2 U891 ( .A1(sh0), .A2(n246), .Z(n662) );
  and2 U892 ( .A1(n125), .A2(n546), .Z(n663) );
  or2 U893 ( .A1(n739), .A2(n740), .Z(n109) );
  and2 U894 ( .A1(inD11), .A2(n918), .Z(n740) );
  and2 U895 ( .A1(inD9), .A2(n70), .Z(n812) );
  and2 U896 ( .A1(n702), .A2(n703), .Z(n408) );
  and2 U897 ( .A1(inD15), .A2(n918), .Z(n757) );
  and2 U898 ( .A1(n114), .A2(n553), .Z(n552) );
  or2 U899 ( .A1(n554), .A2(n555), .Z(n553) );
  or2 U900 ( .A1(n560), .A2(n561), .Z(n554) );
  and2 U901 ( .A1(n62), .A2(n636), .Z(n635) );
  and2 U902 ( .A1(n746), .A2(n96), .Z(n733) );
  or2 U903 ( .A1(n93), .A2(n924), .Z(n922) );
  and2 U904 ( .A1(n114), .A2(n115), .Z(n113) );
  and2 U905 ( .A1(n181), .A2(n180), .Z(n177) );
  and2 U906 ( .A1(n58), .A2(n157), .Z(n156) );
  or2 U907 ( .A1(n223), .A2(n224), .Z(n222) );
  and2 U908 ( .A1(n182), .A2(n225), .Z(n224) );
  and2 U909 ( .A1(n226), .A2(n183), .Z(n223) );
  or2 U910 ( .A1(n358), .A2(n359), .Z(n357) );
  or2 U911 ( .A1(n361), .A2(n362), .Z(n360) );
  or2 U912 ( .A1(n426), .A2(n427), .Z(n425) );
  or2 U913 ( .A1(n808), .A2(n809), .Z(n807) );
  inv1 U914 ( .I(musel2), .ZN(n931) );
  inv1 U915 ( .I(n497), .ZN(n911) );
  and2 U916 ( .A1(n690), .A2(n691), .Z(n689) );
  inv1 U917 ( .I(n419), .ZN(n905) );
  inv1 U918 ( .I(n905), .ZN(n907) );
  inv1 U919 ( .I(n905), .ZN(n906) );
  buf0 U920 ( .I(n83), .Z(n908) );
  or2f U921 ( .A1(n276), .A2(n277), .Z(n228) );
  or2f U922 ( .A1(n940), .A2(n941), .Z(n909) );
  or2f U923 ( .A1(n940), .A2(n941), .Z(n910) );
  inv1f U924 ( .I(n911), .ZN(n912) );
  inv1 U925 ( .I(n911), .ZN(n913) );
  and2f U926 ( .A1(n931), .A2(musel1), .Z(n914) );
  and2f U927 ( .A1(n931), .A2(musel1), .Z(n915) );
  or2f U928 ( .A1(n940), .A2(n941), .Z(n916) );
  or2f U929 ( .A1(n940), .A2(n941), .Z(n917) );
  inv1f U930 ( .I(n939), .ZN(n490) );
  or2 U931 ( .A1(n876), .A2(n877), .Z(n919) );
  and2 U932 ( .A1(n135), .A2(n714), .Z(n690) );
  inv1 U933 ( .I(n494), .ZN(n941) );
  and2 U934 ( .A1(n719), .A2(n494), .Z(n717) );
  and2 U935 ( .A1(n912), .A2(inC9), .Z(n720) );
  and2 U936 ( .A1(n913), .A2(inC3), .Z(n699) );
  and2 U937 ( .A1(n912), .A2(inC2), .Z(n707) );
  or2 U938 ( .A1(n708), .A2(n709), .Z(n653) );
  inv1 U939 ( .I(n711), .ZN(n708) );
  or2 U940 ( .A1(n727), .A2(n728), .Z(n688) );
  inv1 U941 ( .I(n730), .ZN(n727) );
  and2 U942 ( .A1(inB11), .A2(n906), .Z(n739) );
  or2 U943 ( .A1(n119), .A2(n120), .Z(n105) );
  or2 U944 ( .A1(n121), .A2(n122), .Z(n120) );
  or2 U945 ( .A1(n721), .A2(n722), .Z(n135) );
  inv1 U946 ( .I(n724), .ZN(n721) );
  and2 U947 ( .A1(n362), .A2(n361), .Z(n358) );
  inv1 U948 ( .I(n360), .ZN(n359) );
  inv1 U949 ( .I(n653), .ZN(n938) );
  and2 U950 ( .A1(n792), .A2(n494), .Z(n791) );
  and2 U951 ( .A1(n497), .A2(inC1), .Z(n793) );
  and2 U952 ( .A1(n892), .A2(n494), .Z(n891) );
  and2 U953 ( .A1(n497), .A2(inC0), .Z(n893) );
  or2 U954 ( .A1(n732), .A2(n686), .Z(n731) );
  and2 U955 ( .A1(n913), .A2(inC10), .Z(n732) );
  and2 U956 ( .A1(n914), .A2(inA10), .Z(n686) );
  or2 U957 ( .A1(n758), .A2(n759), .Z(n102) );
  and2 U958 ( .A1(n915), .A2(inA3), .Z(n347) );
  and2 U959 ( .A1(n914), .A2(inA2), .Z(n394) );
  and2 U960 ( .A1(n914), .A2(inA1), .Z(n782) );
  and2 U961 ( .A1(n915), .A2(inA0), .Z(n838) );
  inv1 U962 ( .I(n945), .ZN(n947) );
  inv1 U963 ( .I(n581), .ZN(n944) );
  and2 U964 ( .A1(n123), .A2(n661), .Z(n659) );
  or2 U965 ( .A1(n662), .A2(n663), .Z(n661) );
  and2 U966 ( .A1(n546), .A2(n755), .Z(n107) );
  or2 U967 ( .A1(n741), .A2(n98), .Z(n735) );
  and2 U968 ( .A1(sh0), .A2(n742), .Z(n741) );
  or2 U969 ( .A1(n737), .A2(n738), .Z(n736) );
  or2 U970 ( .A1(n119), .A2(n558), .Z(n737) );
  and2 U971 ( .A1(n102), .A2(n902), .Z(n100) );
  or2 U972 ( .A1(n94), .A2(n60), .Z(n924) );
  or2 U973 ( .A1(n715), .A2(n716), .Z(n90) );
  inv1 U974 ( .I(n718), .ZN(n715) );
  or2 U975 ( .A1(n128), .A2(n129), .Z(n127) );
  or2 U976 ( .A1(n132), .A2(n930), .Z(n130) );
  and2 U977 ( .A1(n133), .A2(n902), .Z(n194) );
  and2 U978 ( .A1(n546), .A2(n755), .Z(n930) );
  or2 U979 ( .A1(n180), .A2(n181), .Z(n179) );
  or2 U980 ( .A1(n185), .A2(n158), .Z(n929) );
  and2 U981 ( .A1(n245), .A2(n246), .Z(n244) );
  or2 U982 ( .A1(n236), .A2(n98), .Z(n231) );
  and2 U983 ( .A1(sh0), .A2(n237), .Z(n236) );
  or2 U984 ( .A1(n227), .A2(n228), .Z(n225) );
  inv1 U985 ( .I(n225), .ZN(n183) );
  and2 U986 ( .A1(n245), .A2(n125), .Z(n292) );
  or2 U987 ( .A1(n119), .A2(n281), .Z(n239) );
  or2 U988 ( .A1(n282), .A2(n283), .Z(n281) );
  or2 U989 ( .A1(n285), .A2(n98), .Z(n280) );
  and2 U990 ( .A1(sh0), .A2(n286), .Z(n285) );
  or2 U991 ( .A1(n590), .A2(n591), .Z(n274) );
  inv1 U992 ( .I(n274), .ZN(n227) );
  or2 U993 ( .A1(n119), .A2(n302), .Z(n288) );
  or2 U994 ( .A1(n303), .A2(n304), .Z(n302) );
  and2 U995 ( .A1(sh0), .A2(n306), .Z(n305) );
  inv1 U996 ( .I(n317), .ZN(n276) );
  and2 U997 ( .A1(n245), .A2(n109), .Z(n379) );
  or2 U998 ( .A1(n371), .A2(n98), .Z(n367) );
  and2 U999 ( .A1(sh0), .A2(n372), .Z(n371) );
  or2 U1000 ( .A1(n282), .A2(n373), .Z(n372) );
  or2 U1001 ( .A1(n119), .A2(n368), .Z(n308) );
  or2 U1002 ( .A1(n129), .A2(n369), .Z(n368) );
  inv1 U1003 ( .I(n696), .ZN(n695) );
  or2 U1004 ( .A1(n119), .A2(n414), .Z(n375) );
  or2 U1005 ( .A1(n415), .A2(n416), .Z(n414) );
  or2 U1006 ( .A1(n420), .A2(n98), .Z(n413) );
  and2 U1007 ( .A1(sh0), .A2(n421), .Z(n420) );
  inv1 U1008 ( .I(n704), .ZN(n703) );
  or2 U1009 ( .A1(n119), .A2(n797), .Z(n424) );
  or2 U1010 ( .A1(n798), .A2(n799), .Z(n797) );
  or2 U1011 ( .A1(n802), .A2(n98), .Z(n796) );
  and2 U1012 ( .A1(sh0), .A2(n803), .Z(n802) );
  or2 U1013 ( .A1(n370), .A2(n804), .Z(n803) );
  or2 U1014 ( .A1(n119), .A2(n862), .Z(n806) );
  or2 U1015 ( .A1(n287), .A2(n863), .Z(n862) );
  or2 U1016 ( .A1(n123), .A2(n864), .Z(n863) );
  or2 U1017 ( .A1(n871), .A2(n415), .Z(n870) );
  and2 U1018 ( .A1(sh2), .A2(n851), .Z(n871) );
  or2 U1019 ( .A1(n756), .A2(n757), .Z(n437) );
  and2 U1020 ( .A1(inB15), .A2(n419), .Z(n756) );
  and2 U1021 ( .A1(n114), .A2(n298), .Z(n297) );
  or2 U1022 ( .A1(n299), .A2(n300), .Z(n298) );
  and2 U1023 ( .A1(n308), .A2(n309), .Z(n299) );
  and2 U1024 ( .A1(n301), .A2(n288), .Z(n300) );
  and2 U1025 ( .A1(n114), .A2(n843), .Z(n815) );
  or2 U1026 ( .A1(n844), .A2(n845), .Z(n843) );
  and2 U1027 ( .A1(n846), .A2(n847), .Z(n845) );
  and2 U1028 ( .A1(n861), .A2(n806), .Z(n844) );
  or2 U1029 ( .A1(n549), .A2(n552), .Z(n926) );
  and2 U1030 ( .A1(n652), .A2(n89), .Z(n631) );
  or2 U1031 ( .A1(n664), .A2(n665), .Z(O10) );
  or2 U1032 ( .A1(n666), .A2(n667), .Z(n665) );
  or2 U1033 ( .A1(n54), .A2(n55), .Z(O9) );
  or2 U1034 ( .A1(n56), .A2(n57), .Z(n55) );
  or2 U1035 ( .A1(n93), .A2(n94), .Z(n63) );
  or2 U1036 ( .A1(n112), .A2(n113), .Z(n111) );
  or2 U1037 ( .A1(n153), .A2(n154), .Z(O7) );
  or2 U1038 ( .A1(n184), .A2(n185), .Z(n160) );
  or2 U1039 ( .A1(n199), .A2(n200), .Z(O6) );
  or2 U1040 ( .A1(n201), .A2(n202), .Z(n200) );
  or2 U1041 ( .A1(n248), .A2(n249), .Z(O5) );
  or2 U1042 ( .A1(n250), .A2(n251), .Z(n249) );
  or2 U1043 ( .A1(n334), .A2(n335), .Z(O3) );
  or2 U1044 ( .A1(n336), .A2(n337), .Z(n335) );
  or2 U1045 ( .A1(n381), .A2(n382), .Z(O2) );
  or2 U1046 ( .A1(n383), .A2(n384), .Z(n382) );
  or2 U1047 ( .A1(n760), .A2(n761), .Z(O1) );
  or2 U1048 ( .A1(n762), .A2(n763), .Z(n761) );
  inv1 U1049 ( .I(n456), .ZN(n951) );
  inv1 U1050 ( .I(musel3), .ZN(n900) );
  inv1 U1051 ( .I(n935), .ZN(n483) );
  or2f U1052 ( .A1(n579), .A2(n934), .Z(n935) );
  or2 U1053 ( .A1(n504), .A2(n920), .Z(O13) );
  or2 U1054 ( .A1(n505), .A2(n502), .Z(n920) );
  and2 U1055 ( .A1(n456), .A2(n946), .Z(n925) );
  inv1 U1056 ( .I(musel3), .ZN(n921) );
  and2f U1057 ( .A1(n922), .A2(n923), .Z(n59) );
  or2 U1058 ( .A1(n60), .A2(n62), .Z(n923) );
  and2 U1059 ( .A1(n943), .A2(n89), .Z(n453) );
  or2f U1060 ( .A1(n184), .A2(n929), .Z(n927) );
  and2f U1061 ( .A1(n927), .A2(n928), .Z(n157) );
  or2 U1062 ( .A1(n158), .A2(n62), .Z(n928) );
  and2f U1063 ( .A1(n482), .A2(n89), .Z(n932) );
  or2f U1064 ( .A1(n932), .A2(n933), .Z(O14) );
  or2 U1065 ( .A1(n459), .A2(n462), .Z(n933) );
  and2 U1066 ( .A1(n888), .A2(n889), .Z(n949) );
  and2f U1067 ( .A1(n705), .A2(n909), .Z(n704) );
  or2 U1068 ( .A1(n942), .A2(n455), .Z(n934) );
  or2f U1069 ( .A1(n582), .A2(n947), .Z(n946) );
  or2f U1070 ( .A1(n596), .A2(n597), .Z(n317) );
  and2f U1071 ( .A1(n109), .A2(n902), .Z(n128) );
  and2f U1072 ( .A1(n455), .A2(n950), .Z(n936) );
  or2f U1073 ( .A1(n938), .A2(n277), .Z(n937) );
  inv1f U1074 ( .I(n937), .ZN(n691) );
  inv1 U1075 ( .I(n277), .ZN(n318) );
  and2f U1076 ( .A1(n951), .A2(n943), .Z(n526) );
  and2 U1077 ( .A1(n276), .A2(n318), .Z(n315) );
  and2f U1078 ( .A1(n697), .A2(n917), .Z(n696) );
  inv1f U1079 ( .I(n790), .ZN(n789) );
  or2f U1080 ( .A1(n940), .A2(n941), .Z(n939) );
  inv1f U1081 ( .I(n894), .ZN(n940) );
  inv1 U1082 ( .I(n689), .ZN(n948) );
  inv1 U1083 ( .I(n579), .ZN(n531) );
  and2 U1084 ( .A1(n915), .A2(inA9), .Z(n71) );
  or2 U1085 ( .A1(n952), .A2(n951), .Z(n942) );
  inv1f U1086 ( .I(n946), .ZN(n943) );
  inv1 U1087 ( .I(n530), .ZN(n952) );
  and2 U1088 ( .A1(n598), .A2(n910), .Z(n597) );
  and2 U1089 ( .A1(n723), .A2(n939), .Z(n722) );
  and2 U1090 ( .A1(n710), .A2(n939), .Z(n709) );
  or2f U1091 ( .A1(n579), .A2(n942), .Z(n950) );
  and2 U1092 ( .A1(n530), .A2(n579), .Z(n578) );
  or2 U1093 ( .A1(n917), .A2(n717), .Z(n718) );
  or2 U1094 ( .A1(n916), .A2(n705), .Z(n702) );
  or2 U1095 ( .A1(n917), .A2(n697), .Z(n694) );
  or2 U1096 ( .A1(n939), .A2(n723), .Z(n724) );
  or2 U1097 ( .A1(n939), .A2(n710), .Z(n711) );
  and2 U1098 ( .A1(n729), .A2(n916), .Z(n728) );
  and2 U1099 ( .A1(n717), .A2(n910), .Z(n716) );
  or2 U1100 ( .A1(n909), .A2(n729), .Z(n730) );
  and2 U1101 ( .A1(inB13), .A2(n907), .Z(n744) );
  inv1 U1102 ( .I(opsel2), .ZN(n576) );
  or2 U1103 ( .A1(n571), .A2(n572), .Z(n136) );
  and2 U1104 ( .A1(n575), .A2(n576), .Z(n571) );
  and2 U1105 ( .A1(n62), .A2(n573), .Z(n572) );
  and2 U1106 ( .A1(n574), .A2(opsel2), .Z(n573) );
  or2 U1107 ( .A1(n839), .A2(n840), .Z(n65) );
  and2 U1108 ( .A1(opsel1), .A2(n842), .Z(n839) );
  and2 U1109 ( .A1(opsel0), .A2(n841), .Z(n840) );
  inv1 U1110 ( .I(opsel0), .ZN(n842) );
  or2 U1111 ( .A1(n882), .A2(n92), .Z(n114) );
  and2 U1112 ( .A1(n62), .A2(n58), .Z(n882) );
  and2 U1113 ( .A1(n576), .A2(opsel3), .Z(n58) );
  and2 U1114 ( .A1(n501), .A2(n109), .Z(n657) );
  or2 U1115 ( .A1(n241), .A2(n242), .Z(n240) );
  or2 U1116 ( .A1(n290), .A2(n291), .Z(n289) );
  or2 U1117 ( .A1(n377), .A2(n378), .Z(n376) );
  inv1 U1118 ( .I(sh0), .ZN(n546) );
  and2 U1119 ( .A1(musel1), .A2(musel2), .Z(n828) );
  inv1 U1120 ( .I(sh1), .ZN(n547) );
  and2 U1121 ( .A1(inB7), .A2(n906), .Z(n417) );
  and2 U1122 ( .A1(inB6), .A2(n907), .Z(n800) );
  and2 U1123 ( .A1(inB12), .A2(n419), .Z(n758) );
  and2 U1124 ( .A1(n600), .A2(n494), .Z(n598) );
  or2 U1125 ( .A1(n601), .A2(n324), .Z(n600) );
  and2 U1126 ( .A1(n913), .A2(inC4), .Z(n601) );
  and2 U1127 ( .A1(inB4), .A2(n906), .Z(n852) );
  and2 U1128 ( .A1(inB9), .A2(n906), .Z(n811) );
  and2 U1129 ( .A1(inB3), .A2(n907), .Z(n872) );
  and2 U1130 ( .A1(inB0), .A2(n906), .Z(n874) );
  inv1 U1131 ( .I(sh2), .ZN(n902) );
  and2 U1132 ( .A1(n902), .A2(sh1), .Z(n123) );
  and2 U1133 ( .A1(sh1), .A2(sh2), .Z(n119) );
  and2 U1134 ( .A1(inB2), .A2(n907), .Z(n859) );
  and2 U1135 ( .A1(n546), .A2(sh2), .Z(n245) );
  and2 U1136 ( .A1(n547), .A2(n546), .Z(n243) );
  and2 U1137 ( .A1(n902), .A2(n546), .Z(n108) );
  and2 U1138 ( .A1(inB14), .A2(n907), .Z(n750) );
  and2 U1139 ( .A1(n547), .A2(sh0), .Z(n98) );
  and2 U1140 ( .A1(n574), .A2(n883), .Z(n575) );
  or2 U1141 ( .A1(n435), .A2(n436), .Z(n434) );
  and2 U1142 ( .A1(n62), .A2(n437), .Z(n436) );
  and2 U1143 ( .A1(n65), .A2(n438), .Z(n435) );
  or2 U1144 ( .A1(n439), .A2(n440), .Z(n438) );
  and2 U1145 ( .A1(n455), .A2(n456), .Z(n454) );
  inv1 U1146 ( .I(n457), .ZN(n455) );
  or2 U1147 ( .A1(n498), .A2(n499), .Z(n466) );
  and2 U1148 ( .A1(n501), .A2(n246), .Z(n498) );
  and2 U1149 ( .A1(n500), .A2(n437), .Z(n499) );
  or2 U1150 ( .A1(n464), .A2(n465), .Z(n463) );
  and2 U1151 ( .A1(n65), .A2(n467), .Z(n464) );
  and2 U1152 ( .A1(n62), .A2(n466), .Z(n465) );
  or2 U1153 ( .A1(n468), .A2(n469), .Z(n467) );
  or2 U1154 ( .A1(n538), .A2(n539), .Z(n509) );
  and2 U1155 ( .A1(n501), .A2(n125), .Z(n538) );
  or2 U1156 ( .A1(n540), .A2(n541), .Z(n539) );
  and2 U1157 ( .A1(n548), .A2(n246), .Z(n540) );
  or2 U1158 ( .A1(n507), .A2(n508), .Z(n506) );
  and2 U1159 ( .A1(n510), .A2(n65), .Z(n507) );
  and2 U1160 ( .A1(n62), .A2(n509), .Z(n508) );
  or2 U1161 ( .A1(n511), .A2(n512), .Z(n510) );
  or2 U1162 ( .A1(n618), .A2(n619), .Z(n617) );
  and2 U1163 ( .A1(n614), .A2(n72), .Z(n618) );
  and2 U1164 ( .A1(inC12), .A2(n919), .Z(n619) );
  or2 U1165 ( .A1(n620), .A2(n621), .Z(n616) );
  and2 U1166 ( .A1(inA12), .A2(n75), .Z(n621) );
  and2 U1167 ( .A1(n622), .A2(n623), .Z(n620) );
  and2 U1168 ( .A1(n624), .A2(n625), .Z(n623) );
  or2 U1169 ( .A1(n556), .A2(n557), .Z(n555) );
  and2 U1170 ( .A1(n653), .A2(n948), .Z(n652) );
  or2 U1171 ( .A1(n634), .A2(n635), .Z(n633) );
  and2 U1172 ( .A1(n65), .A2(n637), .Z(n634) );
  and2 U1173 ( .A1(n688), .A2(n948), .Z(n687) );
  and2 U1174 ( .A1(n65), .A2(n672), .Z(n669) );
  and2 U1175 ( .A1(n90), .A2(n948), .Z(n88) );
  and2 U1176 ( .A1(n64), .A2(n65), .Z(n60) );
  and2 U1177 ( .A1(n65), .A2(n161), .Z(n158) );
  and2 U1178 ( .A1(n65), .A2(n207), .Z(n204) );
  or2 U1179 ( .A1(n272), .A2(n273), .Z(n271) );
  and2 U1180 ( .A1(n274), .A2(n228), .Z(n273) );
  and2 U1181 ( .A1(n227), .A2(n275), .Z(n272) );
  inv1 U1182 ( .I(n228), .ZN(n275) );
  and2 U1183 ( .A1(n256), .A2(n65), .Z(n253) );
  and2 U1184 ( .A1(n314), .A2(n136), .Z(n296) );
  or2 U1185 ( .A1(n315), .A2(n316), .Z(n314) );
  and2 U1186 ( .A1(n317), .A2(n277), .Z(n316) );
  or2 U1187 ( .A1(n320), .A2(n321), .Z(n319) );
  or2 U1188 ( .A1(n325), .A2(n326), .Z(n320) );
  or2 U1189 ( .A1(n322), .A2(n323), .Z(n321) );
  and2 U1190 ( .A1(inA4), .A2(n75), .Z(n326) );
  and2 U1191 ( .A1(n65), .A2(n58), .Z(n137) );
  and2 U1192 ( .A1(n65), .A2(n342), .Z(n339) );
  or2 U1193 ( .A1(n405), .A2(n406), .Z(n404) );
  and2 U1194 ( .A1(n363), .A2(n407), .Z(n406) );
  and2 U1195 ( .A1(n408), .A2(n364), .Z(n405) );
  and2 U1196 ( .A1(n65), .A2(n389), .Z(n386) );
  and2 U1197 ( .A1(n575), .A2(opsel2), .Z(n92) );
  or2 U1198 ( .A1(n784), .A2(n785), .Z(n783) );
  and2 U1199 ( .A1(n409), .A2(n787), .Z(n784) );
  inv1 U1200 ( .I(n786), .ZN(n785) );
  or2 U1201 ( .A1(n409), .A2(n787), .Z(n786) );
  and2 U1202 ( .A1(n768), .A2(n65), .Z(n765) );
  and2 U1203 ( .A1(n137), .A2(n817), .Z(n816) );
  or2 U1204 ( .A1(n818), .A2(n819), .Z(n817) );
  or2 U1205 ( .A1(n836), .A2(n837), .Z(n818) );
  or2 U1206 ( .A1(n820), .A2(n821), .Z(n819) );
  or2 U1207 ( .A1(n885), .A2(n886), .Z(n884) );
  and2 U1208 ( .A1(n949), .A2(n490), .Z(n885) );
  inv1 U1209 ( .I(n887), .ZN(n886) );
  or2 U1210 ( .A1(n949), .A2(n490), .Z(n887) );
  inv1 U1211 ( .I(n896), .ZN(n89) );
  or2 U1212 ( .A1(opsel3), .A2(n897), .Z(n896) );
  or2 U1213 ( .A1(n898), .A2(n899), .Z(n897) );
  and2 U1214 ( .A1(opsel2), .A2(n883), .Z(n898) );
  or2 U1215 ( .A1(inC11), .A2(n903), .Z(n646) );
  or2 U1216 ( .A1(inB11), .A2(n908), .Z(n647) );
  or2 U1217 ( .A1(inD11), .A2(n921), .Z(n648) );
  or2 U1218 ( .A1(inA11), .A2(n904), .Z(n645) );
  or2 U1219 ( .A1(inC10), .A2(n903), .Z(n681) );
  or2 U1220 ( .A1(inB10), .A2(n908), .Z(n682) );
  or2 U1221 ( .A1(inD10), .A2(n921), .Z(n683) );
  or2 U1222 ( .A1(inA10), .A2(n904), .Z(n680) );
  or2 U1223 ( .A1(inC9), .A2(n903), .Z(n81) );
  or2 U1224 ( .A1(inB9), .A2(n83), .Z(n82) );
  or2 U1225 ( .A1(inD9), .A2(n921), .Z(n86) );
  or2 U1226 ( .A1(inA9), .A2(n904), .Z(n79) );
  and2 U1227 ( .A1(n496), .A2(inA7), .Z(n166) );
  or2 U1228 ( .A1(inC7), .A2(n903), .Z(n173) );
  or2 U1229 ( .A1(inB7), .A2(n83), .Z(n174) );
  or2 U1230 ( .A1(inD7), .A2(n921), .Z(n175) );
  or2 U1231 ( .A1(inA7), .A2(n904), .Z(n172) );
  and2 U1232 ( .A1(n496), .A2(inA6), .Z(n212) );
  or2 U1233 ( .A1(inC6), .A2(n903), .Z(n219) );
  or2 U1234 ( .A1(inB6), .A2(n908), .Z(n220) );
  or2 U1235 ( .A1(inD6), .A2(n921), .Z(n221) );
  or2 U1236 ( .A1(inA6), .A2(n904), .Z(n218) );
  or2 U1237 ( .A1(inC5), .A2(n903), .Z(n265) );
  or2 U1238 ( .A1(inB5), .A2(n908), .Z(n266) );
  or2 U1239 ( .A1(inD5), .A2(n921), .Z(n267) );
  or2 U1240 ( .A1(inA5), .A2(n904), .Z(n264) );
  or2 U1241 ( .A1(inC3), .A2(n903), .Z(n354) );
  or2 U1242 ( .A1(inB3), .A2(n908), .Z(n355) );
  or2 U1243 ( .A1(inD3), .A2(n921), .Z(n356) );
  or2 U1244 ( .A1(inA3), .A2(n904), .Z(n353) );
  or2 U1245 ( .A1(inC2), .A2(n903), .Z(n401) );
  or2 U1246 ( .A1(inB2), .A2(n908), .Z(n402) );
  or2 U1247 ( .A1(inD2), .A2(n921), .Z(n403) );
  or2 U1248 ( .A1(inA2), .A2(n904), .Z(n400) );
  or2 U1249 ( .A1(inC1), .A2(n903), .Z(n777) );
  or2 U1250 ( .A1(inB1), .A2(n908), .Z(n778) );
  or2 U1251 ( .A1(inD1), .A2(n921), .Z(n779) );
  or2 U1252 ( .A1(inA1), .A2(n904), .Z(n776) );
  and2 U1253 ( .A1(musel3), .A2(n835), .Z(n834) );
  or2 U1254 ( .A1(musel1), .A2(musel2), .Z(n835) );
  or2 U1255 ( .A1(inA15), .A2(n904), .Z(n446) );
  and2 U1256 ( .A1(n447), .A2(n448), .Z(n445) );
  or2 U1257 ( .A1(inB15), .A2(n908), .Z(n448) );
  or2 U1258 ( .A1(inC15), .A2(n903), .Z(n447) );
  and2 U1259 ( .A1(n85), .A2(n449), .Z(n443) );
  or2 U1260 ( .A1(inD15), .A2(n921), .Z(n449) );
  and2 U1261 ( .A1(n536), .A2(n494), .Z(n534) );
  or2 U1262 ( .A1(n537), .A2(n515), .Z(n536) );
  and2 U1263 ( .A1(n913), .A2(inC13), .Z(n537) );
  and2 U1264 ( .A1(n915), .A2(inA14), .Z(n472) );
  or2 U1265 ( .A1(inA14), .A2(n904), .Z(n478) );
  and2 U1266 ( .A1(n479), .A2(n480), .Z(n477) );
  or2 U1267 ( .A1(inB14), .A2(n908), .Z(n480) );
  or2 U1268 ( .A1(inC14), .A2(n903), .Z(n479) );
  and2 U1269 ( .A1(n85), .A2(n481), .Z(n475) );
  or2 U1270 ( .A1(inD14), .A2(n921), .Z(n481) );
  and2 U1271 ( .A1(n493), .A2(n494), .Z(n491) );
  or2 U1272 ( .A1(n495), .A2(n472), .Z(n493) );
  and2 U1273 ( .A1(n912), .A2(inC14), .Z(n495) );
  and2 U1274 ( .A1(sh1), .A2(n546), .Z(n545) );
  and2 U1275 ( .A1(n915), .A2(inA13), .Z(n515) );
  or2 U1276 ( .A1(inA13), .A2(n904), .Z(n521) );
  and2 U1277 ( .A1(n522), .A2(n523), .Z(n520) );
  or2 U1278 ( .A1(inB13), .A2(n908), .Z(n523) );
  or2 U1279 ( .A1(inC13), .A2(n903), .Z(n522) );
  and2 U1280 ( .A1(n85), .A2(n524), .Z(n518) );
  or2 U1281 ( .A1(inD13), .A2(n921), .Z(n524) );
  and2 U1282 ( .A1(n612), .A2(n494), .Z(n610) );
  or2 U1283 ( .A1(n613), .A2(n614), .Z(n612) );
  and2 U1284 ( .A1(n912), .A2(inC12), .Z(n613) );
  and2 U1285 ( .A1(n102), .A2(n547), .Z(n565) );
  or2 U1286 ( .A1(n569), .A2(n102), .Z(n559) );
  or2 U1287 ( .A1(n547), .A2(n546), .Z(n569) );
  and2 U1288 ( .A1(n712), .A2(n494), .Z(n710) );
  or2 U1289 ( .A1(n713), .A2(n651), .Z(n712) );
  and2 U1290 ( .A1(n913), .A2(inC11), .Z(n713) );
  and2 U1291 ( .A1(n915), .A2(inA11), .Z(n651) );
  and2 U1292 ( .A1(inC11), .A2(n919), .Z(n640) );
  and2 U1293 ( .A1(n642), .A2(n643), .Z(n641) );
  and2 U1294 ( .A1(n644), .A2(n645), .Z(n643) );
  and2 U1295 ( .A1(n85), .A2(n648), .Z(n642) );
  and2 U1296 ( .A1(n646), .A2(n647), .Z(n644) );
  and2 U1297 ( .A1(n75), .A2(inA11), .Z(n649) );
  and2 U1298 ( .A1(n731), .A2(n494), .Z(n729) );
  and2 U1299 ( .A1(inC10), .A2(n918), .Z(n675) );
  and2 U1300 ( .A1(n677), .A2(n678), .Z(n676) );
  and2 U1301 ( .A1(n679), .A2(n680), .Z(n678) );
  and2 U1302 ( .A1(n85), .A2(n683), .Z(n677) );
  and2 U1303 ( .A1(n681), .A2(n682), .Z(n679) );
  and2 U1304 ( .A1(n75), .A2(inA10), .Z(n684) );
  or2 U1305 ( .A1(n720), .A2(n71), .Z(n719) );
  and2 U1306 ( .A1(inC9), .A2(n918), .Z(n69) );
  and2 U1307 ( .A1(n71), .A2(n72), .Z(n68) );
  and2 U1308 ( .A1(n76), .A2(n77), .Z(n73) );
  and2 U1309 ( .A1(n78), .A2(n79), .Z(n77) );
  and2 U1310 ( .A1(n85), .A2(n86), .Z(n76) );
  and2 U1311 ( .A1(n81), .A2(n82), .Z(n78) );
  inv1 U1312 ( .I(n496), .ZN(n904) );
  inv1 U1313 ( .I(n828), .ZN(n903) );
  or2 U1314 ( .A1(musel3), .A2(musel1), .Z(n83) );
  and2 U1315 ( .A1(n725), .A2(n494), .Z(n723) );
  or2 U1316 ( .A1(n726), .A2(n143), .Z(n725) );
  and2 U1317 ( .A1(n912), .A2(inC8), .Z(n726) );
  and2 U1318 ( .A1(n587), .A2(n494), .Z(n586) );
  or2 U1319 ( .A1(n588), .A2(n166), .Z(n587) );
  and2 U1320 ( .A1(n913), .A2(inC7), .Z(n588) );
  and2 U1321 ( .A1(inC7), .A2(n919), .Z(n165) );
  and2 U1322 ( .A1(n166), .A2(n72), .Z(n164) );
  and2 U1323 ( .A1(n169), .A2(n170), .Z(n167) );
  and2 U1324 ( .A1(n171), .A2(n172), .Z(n170) );
  and2 U1325 ( .A1(n85), .A2(n175), .Z(n169) );
  and2 U1326 ( .A1(n173), .A2(n174), .Z(n171) );
  and2 U1327 ( .A1(n606), .A2(n494), .Z(n604) );
  or2 U1328 ( .A1(n607), .A2(n212), .Z(n606) );
  and2 U1329 ( .A1(n913), .A2(inC6), .Z(n607) );
  and2 U1330 ( .A1(inC6), .A2(n918), .Z(n211) );
  and2 U1331 ( .A1(n212), .A2(n72), .Z(n210) );
  and2 U1332 ( .A1(n215), .A2(n216), .Z(n213) );
  and2 U1333 ( .A1(n217), .A2(n218), .Z(n216) );
  and2 U1334 ( .A1(n85), .A2(n221), .Z(n215) );
  and2 U1335 ( .A1(n219), .A2(n220), .Z(n217) );
  and2 U1336 ( .A1(n594), .A2(n494), .Z(n592) );
  or2 U1337 ( .A1(n595), .A2(n270), .Z(n594) );
  and2 U1338 ( .A1(n912), .A2(inC5), .Z(n595) );
  and2 U1339 ( .A1(n496), .A2(inA5), .Z(n270) );
  and2 U1340 ( .A1(inC5), .A2(n919), .Z(n259) );
  and2 U1341 ( .A1(n261), .A2(n262), .Z(n260) );
  and2 U1342 ( .A1(n263), .A2(n264), .Z(n262) );
  and2 U1343 ( .A1(n85), .A2(n267), .Z(n261) );
  and2 U1344 ( .A1(n265), .A2(n266), .Z(n263) );
  and2 U1345 ( .A1(inA5), .A2(n75), .Z(n268) );
  and2 U1346 ( .A1(n496), .A2(inA4), .Z(n324) );
  or2 U1347 ( .A1(inC4), .A2(n903), .Z(n331) );
  or2 U1348 ( .A1(inB4), .A2(n908), .Z(n332) );
  or2 U1349 ( .A1(inD4), .A2(n921), .Z(n333) );
  or2 U1350 ( .A1(inA4), .A2(n904), .Z(n330) );
  and2 U1351 ( .A1(inB5), .A2(n906), .Z(n867) );
  and2 U1352 ( .A1(inC3), .A2(n70), .Z(n346) );
  and2 U1353 ( .A1(n347), .A2(n72), .Z(n345) );
  and2 U1354 ( .A1(n350), .A2(n351), .Z(n348) );
  and2 U1355 ( .A1(n352), .A2(n353), .Z(n351) );
  and2 U1356 ( .A1(n85), .A2(n356), .Z(n350) );
  and2 U1357 ( .A1(n354), .A2(n355), .Z(n352) );
  and2 U1358 ( .A1(inB10), .A2(n906), .Z(n752) );
  and2 U1359 ( .A1(inC2), .A2(n919), .Z(n393) );
  and2 U1360 ( .A1(n394), .A2(n72), .Z(n392) );
  and2 U1361 ( .A1(n397), .A2(n398), .Z(n395) );
  and2 U1362 ( .A1(n399), .A2(n400), .Z(n398) );
  and2 U1363 ( .A1(n85), .A2(n403), .Z(n397) );
  and2 U1364 ( .A1(n401), .A2(n402), .Z(n399) );
  inv1 U1365 ( .I(opsel3), .ZN(n574) );
  or2 U1366 ( .A1(n949), .A2(n939), .Z(n410) );
  and2 U1367 ( .A1(inC1), .A2(n918), .Z(n771) );
  and2 U1368 ( .A1(n773), .A2(n774), .Z(n772) );
  and2 U1369 ( .A1(n775), .A2(n776), .Z(n774) );
  and2 U1370 ( .A1(n85), .A2(n779), .Z(n773) );
  and2 U1371 ( .A1(n777), .A2(n778), .Z(n775) );
  and2 U1372 ( .A1(n75), .A2(inA1), .Z(n780) );
  inv1 U1373 ( .I(opsel1), .ZN(n841) );
  and2 U1374 ( .A1(inB1), .A2(n907), .Z(n865) );
  and2 U1375 ( .A1(inB8), .A2(n907), .Z(n857) );
  or2 U1376 ( .A1(inC0), .A2(n903), .Z(n826) );
  or2 U1377 ( .A1(inB0), .A2(n908), .Z(n827) );
  or2 U1378 ( .A1(inD0), .A2(n921), .Z(n829) );
  or2 U1379 ( .A1(inA0), .A2(n904), .Z(n825) );
  and2 U1380 ( .A1(n830), .A2(n831), .Z(n85) );
  and2 U1381 ( .A1(n832), .A2(n833), .Z(n831) );
  or2 U1382 ( .A1(n83), .A2(musel2), .Z(n830) );
  inv1 U1383 ( .I(n834), .ZN(n833) );
  or2 U1384 ( .A1(n497), .A2(n496), .Z(n881) );
  or2 U1385 ( .A1(n441), .A2(n442), .Z(n440) );
  and2 U1386 ( .A1(n443), .A2(n444), .Z(n442) );
  and2 U1387 ( .A1(inC15), .A2(n70), .Z(n441) );
  and2 U1388 ( .A1(n445), .A2(n446), .Z(n444) );
  or2 U1389 ( .A1(n450), .A2(n451), .Z(n439) );
  and2 U1390 ( .A1(n452), .A2(n72), .Z(n451) );
  and2 U1391 ( .A1(n75), .A2(inA15), .Z(n450) );
  or2 U1392 ( .A1(n532), .A2(n533), .Z(n456) );
  and2 U1393 ( .A1(n490), .A2(n535), .Z(n532) );
  and2 U1394 ( .A1(n534), .A2(n939), .Z(n533) );
  inv1 U1395 ( .I(n534), .ZN(n535) );
  or2 U1396 ( .A1(n245), .A2(n658), .Z(n500) );
  or2 U1397 ( .A1(n123), .A2(n98), .Z(n658) );
  or2 U1398 ( .A1(n470), .A2(n471), .Z(n469) );
  and2 U1399 ( .A1(n472), .A2(n72), .Z(n470) );
  and2 U1400 ( .A1(inC14), .A2(n70), .Z(n471) );
  or2 U1401 ( .A1(n473), .A2(n474), .Z(n468) );
  and2 U1402 ( .A1(inA14), .A2(n75), .Z(n474) );
  and2 U1403 ( .A1(n475), .A2(n476), .Z(n473) );
  and2 U1404 ( .A1(n477), .A2(n478), .Z(n476) );
  and2 U1405 ( .A1(n487), .A2(n488), .Z(n457) );
  or2 U1406 ( .A1(n489), .A2(n490), .Z(n488) );
  or2 U1407 ( .A1(n939), .A2(n491), .Z(n487) );
  inv1 U1408 ( .I(n491), .ZN(n489) );
  and2 U1409 ( .A1(n902), .A2(n98), .Z(n548) );
  and2 U1410 ( .A1(n542), .A2(n437), .Z(n541) );
  or2 U1411 ( .A1(n543), .A2(n544), .Z(n542) );
  and2 U1412 ( .A1(sh2), .A2(n547), .Z(n543) );
  or2 U1413 ( .A1(n123), .A2(n545), .Z(n544) );
  or2 U1414 ( .A1(n513), .A2(n514), .Z(n512) );
  and2 U1415 ( .A1(n515), .A2(n72), .Z(n513) );
  and2 U1416 ( .A1(inC13), .A2(n918), .Z(n514) );
  or2 U1417 ( .A1(n516), .A2(n517), .Z(n511) );
  and2 U1418 ( .A1(inA13), .A2(n75), .Z(n517) );
  and2 U1419 ( .A1(n518), .A2(n519), .Z(n516) );
  and2 U1420 ( .A1(n520), .A2(n521), .Z(n519) );
  and2 U1421 ( .A1(n914), .A2(inA12), .Z(n614) );
  or2 U1422 ( .A1(inA12), .A2(n904), .Z(n625) );
  and2 U1423 ( .A1(n626), .A2(n627), .Z(n624) );
  or2 U1424 ( .A1(inB12), .A2(n908), .Z(n627) );
  or2 U1425 ( .A1(inC12), .A2(n903), .Z(n626) );
  and2 U1426 ( .A1(n85), .A2(n628), .Z(n622) );
  or2 U1427 ( .A1(inD12), .A2(n921), .Z(n628) );
  or2 U1428 ( .A1(n608), .A2(n609), .Z(n530) );
  and2 U1429 ( .A1(n490), .A2(n611), .Z(n608) );
  and2 U1430 ( .A1(n610), .A2(n939), .Z(n609) );
  inv1 U1431 ( .I(n610), .ZN(n611) );
  and2 U1432 ( .A1(sh0), .A2(n566), .Z(n560) );
  or2 U1433 ( .A1(n567), .A2(n568), .Z(n566) );
  and2 U1434 ( .A1(n123), .A2(n437), .Z(n568) );
  and2 U1435 ( .A1(n119), .A2(n559), .Z(n567) );
  or2 U1436 ( .A1(n562), .A2(n563), .Z(n561) );
  and2 U1437 ( .A1(n564), .A2(n123), .Z(n563) );
  and2 U1438 ( .A1(n565), .A2(n108), .Z(n562) );
  and2 U1439 ( .A1(n246), .A2(n546), .Z(n564) );
  and2 U1440 ( .A1(n558), .A2(n559), .Z(n557) );
  and2 U1441 ( .A1(n548), .A2(n125), .Z(n556) );
  inv1 U1442 ( .I(n500), .ZN(n501) );
  and2 U1443 ( .A1(n548), .A2(n102), .Z(n660) );
  and2 U1444 ( .A1(n558), .A2(n569), .Z(n656) );
  or2 U1445 ( .A1(n638), .A2(n639), .Z(n637) );
  or2 U1446 ( .A1(n649), .A2(n650), .Z(n638) );
  or2 U1447 ( .A1(n640), .A2(n641), .Z(n639) );
  and2 U1448 ( .A1(n651), .A2(n72), .Z(n650) );
  or2 U1449 ( .A1(n123), .A2(n128), .Z(n738) );
  and2 U1450 ( .A1(n108), .A2(n102), .Z(n754) );
  or2 U1451 ( .A1(n673), .A2(n674), .Z(n672) );
  or2 U1452 ( .A1(n684), .A2(n685), .Z(n673) );
  or2 U1453 ( .A1(n675), .A2(n676), .Z(n674) );
  and2 U1454 ( .A1(n686), .A2(n72), .Z(n685) );
  and2 U1455 ( .A1(n108), .A2(n109), .Z(n106) );
  or2 U1456 ( .A1(n66), .A2(n67), .Z(n64) );
  or2 U1457 ( .A1(n73), .A2(n74), .Z(n66) );
  or2 U1458 ( .A1(n68), .A2(n69), .Z(n67) );
  and2 U1459 ( .A1(n75), .A2(inA9), .Z(n74) );
  and2 U1460 ( .A1(n914), .A2(inA8), .Z(n143) );
  and2 U1461 ( .A1(n879), .A2(n931), .Z(n878) );
  or2 U1462 ( .A1(inA8), .A2(n904), .Z(n149) );
  and2 U1463 ( .A1(n150), .A2(n151), .Z(n148) );
  or2 U1464 ( .A1(inB8), .A2(n908), .Z(n151) );
  or2 U1465 ( .A1(inC8), .A2(n903), .Z(n150) );
  and2 U1466 ( .A1(n85), .A2(n152), .Z(n146) );
  or2 U1467 ( .A1(inD8), .A2(n921), .Z(n152) );
  and2 U1468 ( .A1(n108), .A2(n133), .Z(n132) );
  or2 U1469 ( .A1(n126), .A2(n98), .Z(n118) );
  and2 U1470 ( .A1(sh0), .A2(n127), .Z(n126) );
  and2 U1471 ( .A1(n108), .A2(n198), .Z(n197) );
  and2 U1472 ( .A1(n583), .A2(n584), .Z(n180) );
  or2 U1473 ( .A1(n585), .A2(n490), .Z(n584) );
  or2 U1474 ( .A1(n939), .A2(n586), .Z(n583) );
  inv1 U1475 ( .I(n586), .ZN(n585) );
  or2 U1476 ( .A1(n162), .A2(n163), .Z(n161) );
  or2 U1477 ( .A1(n167), .A2(n168), .Z(n162) );
  or2 U1478 ( .A1(n164), .A2(n165), .Z(n163) );
  and2 U1479 ( .A1(inA7), .A2(n75), .Z(n168) );
  or2 U1480 ( .A1(n243), .A2(n244), .Z(n242) );
  and2 U1481 ( .A1(n108), .A2(n247), .Z(n241) );
  and2 U1482 ( .A1(sh2), .A2(n109), .Z(n233) );
  or2 U1483 ( .A1(n602), .A2(n603), .Z(n182) );
  and2 U1484 ( .A1(n490), .A2(n605), .Z(n602) );
  and2 U1485 ( .A1(n604), .A2(n939), .Z(n603) );
  inv1 U1486 ( .I(n604), .ZN(n605) );
  inv1 U1487 ( .I(n182), .ZN(n226) );
  or2 U1488 ( .A1(n208), .A2(n209), .Z(n207) );
  or2 U1489 ( .A1(n213), .A2(n214), .Z(n208) );
  or2 U1490 ( .A1(n210), .A2(n211), .Z(n209) );
  and2 U1491 ( .A1(inA6), .A2(n75), .Z(n214) );
  or2 U1492 ( .A1(n243), .A2(n292), .Z(n291) );
  and2 U1493 ( .A1(n108), .A2(n293), .Z(n290) );
  and2 U1494 ( .A1(n490), .A2(n593), .Z(n590) );
  and2 U1495 ( .A1(n592), .A2(n939), .Z(n591) );
  inv1 U1496 ( .I(n592), .ZN(n593) );
  or2 U1497 ( .A1(n257), .A2(n258), .Z(n256) );
  or2 U1498 ( .A1(n268), .A2(n269), .Z(n257) );
  or2 U1499 ( .A1(n259), .A2(n260), .Z(n258) );
  and2 U1500 ( .A1(n270), .A2(n72), .Z(n269) );
  or2 U1501 ( .A1(n305), .A2(n98), .Z(n301) );
  or2 U1502 ( .A1(n235), .A2(n307), .Z(n306) );
  or2 U1503 ( .A1(n310), .A2(n311), .Z(n309) );
  and2 U1504 ( .A1(n108), .A2(n313), .Z(n310) );
  or2 U1505 ( .A1(n243), .A2(n312), .Z(n311) );
  and2 U1506 ( .A1(n245), .A2(n102), .Z(n312) );
  and2 U1507 ( .A1(n490), .A2(n599), .Z(n596) );
  inv1 U1508 ( .I(n598), .ZN(n599) );
  and2 U1509 ( .A1(n912), .A2(n72), .Z(n75) );
  and2 U1510 ( .A1(inC4), .A2(n918), .Z(n323) );
  and2 U1511 ( .A1(n324), .A2(n72), .Z(n322) );
  and2 U1512 ( .A1(n327), .A2(n328), .Z(n325) );
  and2 U1513 ( .A1(n329), .A2(n330), .Z(n328) );
  and2 U1514 ( .A1(n85), .A2(n333), .Z(n327) );
  and2 U1515 ( .A1(n331), .A2(n332), .Z(n329) );
  or2 U1516 ( .A1(n243), .A2(n379), .Z(n378) );
  and2 U1517 ( .A1(n108), .A2(n380), .Z(n377) );
  and2 U1518 ( .A1(n363), .A2(n364), .Z(n362) );
  or2 U1519 ( .A1(n343), .A2(n344), .Z(n342) );
  or2 U1520 ( .A1(n348), .A2(n349), .Z(n343) );
  or2 U1521 ( .A1(n345), .A2(n346), .Z(n344) );
  and2 U1522 ( .A1(n75), .A2(inA3), .Z(n349) );
  or2 U1523 ( .A1(n243), .A2(n428), .Z(n427) );
  and2 U1524 ( .A1(n245), .A2(n133), .Z(n428) );
  and2 U1525 ( .A1(n108), .A2(n429), .Z(n426) );
  or2 U1526 ( .A1(n409), .A2(n410), .Z(n407) );
  inv1 U1527 ( .I(n407), .ZN(n364) );
  inv1 U1528 ( .I(n408), .ZN(n363) );
  or2 U1529 ( .A1(n390), .A2(n391), .Z(n389) );
  or2 U1530 ( .A1(n395), .A2(n396), .Z(n390) );
  or2 U1531 ( .A1(n392), .A2(n393), .Z(n391) );
  and2 U1532 ( .A1(n75), .A2(inA2), .Z(n396) );
  or2 U1533 ( .A1(n243), .A2(n810), .Z(n809) );
  and2 U1534 ( .A1(n245), .A2(n198), .Z(n810) );
  and2 U1535 ( .A1(n108), .A2(n374), .Z(n808) );
  and2 U1536 ( .A1(n423), .A2(n902), .Z(n798) );
  inv1 U1537 ( .I(n410), .ZN(n787) );
  inv1 U1538 ( .I(n883), .ZN(n62) );
  or2 U1539 ( .A1(n769), .A2(n770), .Z(n768) );
  or2 U1540 ( .A1(n780), .A2(n781), .Z(n769) );
  or2 U1541 ( .A1(n771), .A2(n772), .Z(n770) );
  and2 U1542 ( .A1(n782), .A2(n72), .Z(n781) );
  or2 U1543 ( .A1(n869), .A2(n98), .Z(n861) );
  and2 U1544 ( .A1(sh0), .A2(n870), .Z(n869) );
  or2 U1545 ( .A1(n848), .A2(n849), .Z(n847) );
  or2 U1546 ( .A1(n123), .A2(n119), .Z(n848) );
  or2 U1547 ( .A1(n307), .A2(n850), .Z(n849) );
  and2 U1548 ( .A1(n851), .A2(n902), .Z(n850) );
  or2 U1549 ( .A1(n854), .A2(n855), .Z(n846) );
  and2 U1550 ( .A1(n108), .A2(n423), .Z(n854) );
  or2 U1551 ( .A1(n243), .A2(n856), .Z(n855) );
  and2 U1552 ( .A1(n245), .A2(n247), .Z(n856) );
  and2 U1553 ( .A1(inC0), .A2(n70), .Z(n820) );
  and2 U1554 ( .A1(n822), .A2(n823), .Z(n821) );
  and2 U1555 ( .A1(n824), .A2(n825), .Z(n823) );
  and2 U1556 ( .A1(n85), .A2(n829), .Z(n822) );
  and2 U1557 ( .A1(n826), .A2(n827), .Z(n824) );
  and2 U1558 ( .A1(n75), .A2(inA0), .Z(n836) );
  and2 U1559 ( .A1(n838), .A2(n72), .Z(n837) );
  or2 U1560 ( .A1(opsel0), .A2(opsel1), .Z(n883) );
  and2 U1561 ( .A1(n62), .A2(n576), .Z(n899) );
  or2 U1562 ( .A1(n141), .A2(n142), .Z(n140) );
  and2 U1563 ( .A1(n143), .A2(n72), .Z(n141) );
  and2 U1564 ( .A1(inC8), .A2(n70), .Z(n142) );
  or2 U1565 ( .A1(n144), .A2(n145), .Z(n139) );
  and2 U1566 ( .A1(n75), .A2(inA8), .Z(n145) );
  and2 U1567 ( .A1(n146), .A2(n147), .Z(n144) );
  and2 U1568 ( .A1(n148), .A2(n149), .Z(n147) );
  or2 U1569 ( .A1(n116), .A2(n117), .Z(n115) );
  and2 U1570 ( .A1(n118), .A2(n105), .Z(n117) );
  and2 U1571 ( .A1(n130), .A2(n131), .Z(n116) );
  and2 U1572 ( .A1(n134), .A2(n135), .Z(n112) );
  and2 U1573 ( .A1(n136), .A2(n948), .Z(n134) );
  and2 U1574 ( .A1(n92), .A2(n437), .Z(n430) );
  and2 U1575 ( .A1(n58), .A2(n434), .Z(n433) );
  and2 U1576 ( .A1(n92), .A2(n466), .Z(n459) );
  and2 U1577 ( .A1(n58), .A2(n463), .Z(n462) );
  and2 U1578 ( .A1(n92), .A2(n509), .Z(n502) );
  and2 U1579 ( .A1(n58), .A2(n506), .Z(n505) );
  and2 U1580 ( .A1(n137), .A2(n615), .Z(n549) );
  or2 U1581 ( .A1(n616), .A2(n617), .Z(n615) );
  or2 U1582 ( .A1(n629), .A2(n630), .Z(O11) );
  and2 U1583 ( .A1(n92), .A2(n636), .Z(n629) );
  or2 U1584 ( .A1(n631), .A2(n632), .Z(n630) );
  and2 U1585 ( .A1(n92), .A2(n671), .Z(n664) );
  and2 U1586 ( .A1(n687), .A2(n89), .Z(n666) );
  and2 U1587 ( .A1(n92), .A2(n63), .Z(n54) );
  and2 U1588 ( .A1(n88), .A2(n89), .Z(n56) );
  or2 U1589 ( .A1(n110), .A2(n111), .Z(O8) );
  and2 U1590 ( .A1(n137), .A2(n138), .Z(n110) );
  or2 U1591 ( .A1(n139), .A2(n140), .Z(n138) );
  and2 U1592 ( .A1(n92), .A2(n160), .Z(n153) );
  and2 U1593 ( .A1(n92), .A2(n206), .Z(n199) );
  and2 U1594 ( .A1(n89), .A2(n222), .Z(n201) );
  and2 U1595 ( .A1(n92), .A2(n255), .Z(n248) );
  and2 U1596 ( .A1(n89), .A2(n271), .Z(n250) );
  and2 U1597 ( .A1(n137), .A2(n319), .Z(n294) );
  or2 U1598 ( .A1(n296), .A2(n297), .Z(n295) );
  and2 U1599 ( .A1(n92), .A2(n341), .Z(n334) );
  and2 U1600 ( .A1(n89), .A2(n357), .Z(n336) );
  and2 U1601 ( .A1(n92), .A2(n388), .Z(n381) );
  and2 U1602 ( .A1(n89), .A2(n404), .Z(n383) );
  and2 U1603 ( .A1(n92), .A2(n767), .Z(n760) );
  and2 U1604 ( .A1(n89), .A2(n783), .Z(n762) );
  and2 U1605 ( .A1(n89), .A2(n884), .Z(n813) );
  or2 U1606 ( .A1(n815), .A2(n816), .Z(n814) );
  or2 U1607 ( .A1(n294), .A2(n295), .Z(O4) );
  or2 U1608 ( .A1(n813), .A2(n814), .Z(O0) );
endmodule

